VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO solo_squash_caravel_gf180
  CLASS BLOCK ;
  FOREIGN solo_squash_caravel_gf180 ;
  ORIGIN 0.000 0.000 ;
  SIZE 209.505 BY 227.425 ;
  PIN blue
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 73.920 209.505 74.480 ;
    END
  END blue
  PIN debug_design_reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 67.200 209.505 67.760 ;
    END
  END debug_design_reset
  PIN debug_gpio_ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 10.080 209.505 10.640 ;
    END
  END debug_gpio_ready
  PIN down_key_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END down_key_n
  PIN ext_reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 131.040 209.505 131.600 ;
    END
  END ext_reset_n
  PIN gpio_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 13.440 209.505 14.000 ;
    END
  END gpio_ready
  PIN green
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 104.160 209.505 104.720 ;
    END
  END green
  PIN hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 100.800 209.505 101.360 ;
    END
  END hsync
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 218.400 209.505 218.960 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 4.000 17.360 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 201.600 209.505 202.160 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 77.280 209.505 77.840 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 87.360 209.505 87.920 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 90.720 209.505 91.280 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 84.000 209.505 84.560 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 94.080 209.505 94.640 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 80.640 209.505 81.200 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 16.800 209.505 17.360 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 20.160 209.505 20.720 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 63.840 209.505 64.400 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 215.040 209.505 215.600 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 40.320 209.505 40.880 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 204.960 209.505 205.520 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 36.960 209.505 37.520 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 223.425 40.880 227.425 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.800 4.000 185.360 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 198.240 209.505 198.800 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 211.680 209.505 212.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 26.880 209.505 27.440 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 191.520 209.505 192.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 208.320 209.505 208.880 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 194.880 209.505 195.440 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 188.160 209.505 188.720 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 223.425 178.640 227.425 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 23.520 209.505 24.080 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 30.240 209.505 30.800 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 33.600 209.505 34.160 ;
    END
  END io_oeb[9]
  PIN new_game_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END new_game_n
  PIN pause_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END pause_n
  PIN red
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 97.440 209.505 98.000 ;
    END
  END red
  PIN speaker
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END speaker
  PIN up_key_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END up_key_n
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 211.980 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 211.980 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 211.980 ;
    END
  END vss
  PIN vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END vsync
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 205.505 134.400 209.505 134.960 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 202.720 211.980 ;
      LAYER Metal2 ;
        RECT 8.540 223.125 40.020 223.425 ;
        RECT 41.180 223.125 177.780 223.425 ;
        RECT 178.940 223.125 202.020 223.425 ;
        RECT 8.540 4.300 202.020 223.125 ;
        RECT 8.540 4.000 50.100 4.300 ;
        RECT 51.260 4.000 53.460 4.300 ;
        RECT 54.620 4.000 97.140 4.300 ;
        RECT 98.300 4.000 100.500 4.300 ;
        RECT 101.660 4.000 164.340 4.300 ;
        RECT 165.500 4.000 202.020 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 218.100 205.205 218.820 ;
        RECT 4.000 215.900 205.505 218.100 ;
        RECT 4.000 214.740 205.205 215.900 ;
        RECT 4.000 212.540 205.505 214.740 ;
        RECT 4.000 211.380 205.205 212.540 ;
        RECT 4.000 209.180 205.505 211.380 ;
        RECT 4.000 208.020 205.205 209.180 ;
        RECT 4.000 205.820 205.505 208.020 ;
        RECT 4.300 204.660 205.205 205.820 ;
        RECT 4.000 202.460 205.505 204.660 ;
        RECT 4.300 201.300 205.205 202.460 ;
        RECT 4.000 199.100 205.505 201.300 ;
        RECT 4.000 197.940 205.205 199.100 ;
        RECT 4.000 195.740 205.505 197.940 ;
        RECT 4.000 194.580 205.205 195.740 ;
        RECT 4.000 192.380 205.505 194.580 ;
        RECT 4.000 191.220 205.205 192.380 ;
        RECT 4.000 189.020 205.505 191.220 ;
        RECT 4.300 187.860 205.205 189.020 ;
        RECT 4.000 185.660 205.505 187.860 ;
        RECT 4.300 184.500 205.505 185.660 ;
        RECT 4.000 135.260 205.505 184.500 ;
        RECT 4.000 134.100 205.205 135.260 ;
        RECT 4.000 131.900 205.505 134.100 ;
        RECT 4.000 130.740 205.205 131.900 ;
        RECT 4.000 125.180 205.505 130.740 ;
        RECT 4.300 124.020 205.505 125.180 ;
        RECT 4.000 121.820 205.505 124.020 ;
        RECT 4.300 120.660 205.505 121.820 ;
        RECT 4.000 105.020 205.505 120.660 ;
        RECT 4.000 103.860 205.205 105.020 ;
        RECT 4.000 101.660 205.505 103.860 ;
        RECT 4.300 100.500 205.205 101.660 ;
        RECT 4.000 98.300 205.505 100.500 ;
        RECT 4.300 97.140 205.205 98.300 ;
        RECT 4.000 94.940 205.505 97.140 ;
        RECT 4.000 93.780 205.205 94.940 ;
        RECT 4.000 91.580 205.505 93.780 ;
        RECT 4.000 90.420 205.205 91.580 ;
        RECT 4.000 88.220 205.505 90.420 ;
        RECT 4.000 87.060 205.205 88.220 ;
        RECT 4.000 84.860 205.505 87.060 ;
        RECT 4.000 83.700 205.205 84.860 ;
        RECT 4.000 81.500 205.505 83.700 ;
        RECT 4.000 80.340 205.205 81.500 ;
        RECT 4.000 78.140 205.505 80.340 ;
        RECT 4.000 76.980 205.205 78.140 ;
        RECT 4.000 74.780 205.505 76.980 ;
        RECT 4.000 73.620 205.205 74.780 ;
        RECT 4.000 68.060 205.505 73.620 ;
        RECT 4.000 66.900 205.205 68.060 ;
        RECT 4.000 64.700 205.505 66.900 ;
        RECT 4.000 63.540 205.205 64.700 ;
        RECT 4.000 41.180 205.505 63.540 ;
        RECT 4.000 40.020 205.205 41.180 ;
        RECT 4.000 37.820 205.505 40.020 ;
        RECT 4.000 36.660 205.205 37.820 ;
        RECT 4.000 34.460 205.505 36.660 ;
        RECT 4.000 33.300 205.205 34.460 ;
        RECT 4.000 31.100 205.505 33.300 ;
        RECT 4.300 29.940 205.205 31.100 ;
        RECT 4.000 27.740 205.505 29.940 ;
        RECT 4.300 26.580 205.205 27.740 ;
        RECT 4.000 24.380 205.505 26.580 ;
        RECT 4.300 23.220 205.205 24.380 ;
        RECT 4.000 21.020 205.505 23.220 ;
        RECT 4.300 19.860 205.205 21.020 ;
        RECT 4.000 17.660 205.505 19.860 ;
        RECT 4.300 16.500 205.205 17.660 ;
        RECT 4.000 14.300 205.505 16.500 ;
        RECT 4.000 13.140 205.205 14.300 ;
        RECT 4.000 10.940 205.505 13.140 ;
        RECT 4.000 10.220 205.205 10.940 ;
      LAYER Metal4 ;
        RECT 21.420 17.450 21.940 176.870 ;
        RECT 24.140 17.450 98.740 176.870 ;
        RECT 100.940 17.450 172.900 176.870 ;
  END
END solo_squash_caravel_gf180
END LIBRARY


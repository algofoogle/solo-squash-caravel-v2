magic
tech gf180mcuD
magscale 1 10
timestamp 1701082017
<< metal1 >>
rect 1344 42362 40544 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 40544 42362
rect 1344 42276 40544 42310
rect 8318 42194 8370 42206
rect 8318 42130 8370 42142
rect 35982 42194 36034 42206
rect 35982 42130 36034 42142
rect 38782 42194 38834 42206
rect 38782 42130 38834 42142
rect 40126 42194 40178 42206
rect 40126 42130 40178 42142
rect 39230 42082 39282 42094
rect 39230 42018 39282 42030
rect 1344 41578 40544 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 40544 41578
rect 1344 41492 40544 41526
rect 39678 41074 39730 41086
rect 39678 41010 39730 41022
rect 1710 40962 1762 40974
rect 1710 40898 1762 40910
rect 29374 40962 29426 40974
rect 29374 40898 29426 40910
rect 30382 40962 30434 40974
rect 30382 40898 30434 40910
rect 30830 40962 30882 40974
rect 30830 40898 30882 40910
rect 40126 40962 40178 40974
rect 40126 40898 40178 40910
rect 1344 40794 40544 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 40544 40794
rect 1344 40708 40544 40742
rect 40126 40514 40178 40526
rect 40126 40450 40178 40462
rect 29150 40402 29202 40414
rect 25890 40350 25902 40402
rect 25954 40350 25966 40402
rect 29586 40350 29598 40402
rect 29650 40350 29662 40402
rect 29150 40338 29202 40350
rect 26562 40238 26574 40290
rect 26626 40238 26638 40290
rect 28690 40238 28702 40290
rect 28754 40238 28766 40290
rect 30370 40238 30382 40290
rect 30434 40238 30446 40290
rect 32498 40238 32510 40290
rect 32562 40238 32574 40290
rect 1344 40010 40544 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 40544 40010
rect 1344 39924 40544 39958
rect 27246 39842 27298 39854
rect 27246 39778 27298 39790
rect 31166 39730 31218 39742
rect 26338 39678 26350 39730
rect 26402 39678 26414 39730
rect 31166 39666 31218 39678
rect 31838 39730 31890 39742
rect 31838 39666 31890 39678
rect 31950 39730 32002 39742
rect 31950 39666 32002 39678
rect 23538 39566 23550 39618
rect 23602 39566 23614 39618
rect 29362 39566 29374 39618
rect 29426 39566 29438 39618
rect 30818 39566 30830 39618
rect 30882 39566 30894 39618
rect 32722 39566 32734 39618
rect 32786 39566 32798 39618
rect 27358 39506 27410 39518
rect 24210 39454 24222 39506
rect 24274 39454 24286 39506
rect 27358 39442 27410 39454
rect 27582 39506 27634 39518
rect 27582 39442 27634 39454
rect 31502 39506 31554 39518
rect 31502 39442 31554 39454
rect 32062 39506 32114 39518
rect 32062 39442 32114 39454
rect 26798 39394 26850 39406
rect 29934 39394 29986 39406
rect 29138 39342 29150 39394
rect 29202 39342 29214 39394
rect 26798 39330 26850 39342
rect 29934 39330 29986 39342
rect 30046 39394 30098 39406
rect 30046 39330 30098 39342
rect 30158 39394 30210 39406
rect 30158 39330 30210 39342
rect 30382 39394 30434 39406
rect 30382 39330 30434 39342
rect 31054 39394 31106 39406
rect 31054 39330 31106 39342
rect 31278 39394 31330 39406
rect 40126 39394 40178 39406
rect 32498 39342 32510 39394
rect 32562 39342 32574 39394
rect 31278 39330 31330 39342
rect 40126 39330 40178 39342
rect 1344 39226 40544 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 40544 39226
rect 1344 39140 40544 39174
rect 25342 39058 25394 39070
rect 29810 39006 29822 39058
rect 29874 39006 29886 39058
rect 25342 38994 25394 39006
rect 33070 38946 33122 38958
rect 31378 38894 31390 38946
rect 31442 38894 31454 38946
rect 32050 38894 32062 38946
rect 32114 38894 32126 38946
rect 33070 38882 33122 38894
rect 33294 38946 33346 38958
rect 33294 38882 33346 38894
rect 40126 38946 40178 38958
rect 40126 38882 40178 38894
rect 32398 38834 32450 38846
rect 11330 38782 11342 38834
rect 11394 38782 11406 38834
rect 25554 38782 25566 38834
rect 25618 38782 25630 38834
rect 28242 38782 28254 38834
rect 28306 38782 28318 38834
rect 30034 38782 30046 38834
rect 30098 38782 30110 38834
rect 30930 38782 30942 38834
rect 30994 38782 31006 38834
rect 32398 38770 32450 38782
rect 25230 38722 25282 38734
rect 28814 38722 28866 38734
rect 12002 38670 12014 38722
rect 12066 38670 12078 38722
rect 14130 38670 14142 38722
rect 14194 38670 14206 38722
rect 27906 38670 27918 38722
rect 27970 38670 27982 38722
rect 25230 38658 25282 38670
rect 28814 38658 28866 38670
rect 33182 38722 33234 38734
rect 33182 38658 33234 38670
rect 1344 38442 40544 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40544 38442
rect 1344 38356 40544 38390
rect 12350 38274 12402 38286
rect 12350 38210 12402 38222
rect 31502 38274 31554 38286
rect 31502 38210 31554 38222
rect 31726 38274 31778 38286
rect 31726 38210 31778 38222
rect 21534 38162 21586 38174
rect 30158 38162 30210 38174
rect 14242 38110 14254 38162
rect 14306 38110 14318 38162
rect 16258 38110 16270 38162
rect 16322 38110 16334 38162
rect 25106 38110 25118 38162
rect 25170 38110 25182 38162
rect 28018 38110 28030 38162
rect 28082 38110 28094 38162
rect 29362 38110 29374 38162
rect 29426 38110 29438 38162
rect 21534 38098 21586 38110
rect 30158 38098 30210 38110
rect 26574 38050 26626 38062
rect 28366 38050 28418 38062
rect 31166 38050 31218 38062
rect 14130 37998 14142 38050
rect 14194 37998 14206 38050
rect 19170 37998 19182 38050
rect 19234 37998 19246 38050
rect 25330 37998 25342 38050
rect 25394 37998 25406 38050
rect 26114 37998 26126 38050
rect 26178 37998 26190 38050
rect 27906 37998 27918 38050
rect 27970 37998 27982 38050
rect 29698 37998 29710 38050
rect 29762 37998 29774 38050
rect 26574 37986 26626 37998
rect 28366 37986 28418 37998
rect 31166 37986 31218 37998
rect 12686 37938 12738 37950
rect 12686 37874 12738 37886
rect 13470 37938 13522 37950
rect 13470 37874 13522 37886
rect 15486 37938 15538 37950
rect 21422 37938 21474 37950
rect 18386 37886 18398 37938
rect 18450 37886 18462 37938
rect 15486 37874 15538 37886
rect 21422 37874 21474 37886
rect 21646 37938 21698 37950
rect 21646 37874 21698 37886
rect 24670 37938 24722 37950
rect 24670 37874 24722 37886
rect 25118 37938 25170 37950
rect 25118 37874 25170 37886
rect 26686 37938 26738 37950
rect 26686 37874 26738 37886
rect 27358 37938 27410 37950
rect 27358 37874 27410 37886
rect 28590 37938 28642 37950
rect 28590 37874 28642 37886
rect 30494 37938 30546 37950
rect 30494 37874 30546 37886
rect 30942 37938 30994 37950
rect 30942 37874 30994 37886
rect 12462 37826 12514 37838
rect 12462 37762 12514 37774
rect 14814 37826 14866 37838
rect 15598 37826 15650 37838
rect 15138 37774 15150 37826
rect 15202 37774 15214 37826
rect 14814 37762 14866 37774
rect 15598 37762 15650 37774
rect 15822 37826 15874 37838
rect 15822 37762 15874 37774
rect 19630 37826 19682 37838
rect 19630 37762 19682 37774
rect 24894 37826 24946 37838
rect 24894 37762 24946 37774
rect 28142 37826 28194 37838
rect 28142 37762 28194 37774
rect 30606 37826 30658 37838
rect 30606 37762 30658 37774
rect 31838 37826 31890 37838
rect 31838 37762 31890 37774
rect 32174 37826 32226 37838
rect 40126 37826 40178 37838
rect 32498 37774 32510 37826
rect 32562 37774 32574 37826
rect 32174 37762 32226 37774
rect 40126 37762 40178 37774
rect 1344 37658 40544 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40544 37658
rect 1344 37572 40544 37606
rect 9662 37490 9714 37502
rect 9662 37426 9714 37438
rect 17614 37490 17666 37502
rect 28030 37490 28082 37502
rect 23202 37438 23214 37490
rect 23266 37438 23278 37490
rect 27458 37438 27470 37490
rect 27522 37438 27534 37490
rect 17614 37426 17666 37438
rect 28030 37426 28082 37438
rect 30606 37490 30658 37502
rect 30606 37426 30658 37438
rect 31278 37490 31330 37502
rect 31278 37426 31330 37438
rect 1710 37378 1762 37390
rect 1710 37314 1762 37326
rect 16718 37378 16770 37390
rect 16718 37314 16770 37326
rect 17390 37378 17442 37390
rect 30382 37378 30434 37390
rect 40126 37378 40178 37390
rect 21746 37326 21758 37378
rect 21810 37326 21822 37378
rect 26562 37326 26574 37378
rect 26626 37326 26638 37378
rect 32050 37326 32062 37378
rect 32114 37326 32126 37378
rect 17390 37314 17442 37326
rect 30382 37314 30434 37326
rect 40126 37314 40178 37326
rect 16158 37266 16210 37278
rect 13458 37214 13470 37266
rect 13522 37214 13534 37266
rect 15474 37214 15486 37266
rect 15538 37214 15550 37266
rect 16158 37202 16210 37214
rect 16382 37266 16434 37278
rect 22878 37266 22930 37278
rect 30270 37266 30322 37278
rect 17826 37214 17838 37266
rect 17890 37214 17902 37266
rect 22530 37214 22542 37266
rect 22594 37214 22606 37266
rect 26450 37214 26462 37266
rect 26514 37214 26526 37266
rect 27346 37214 27358 37266
rect 27410 37214 27422 37266
rect 16382 37202 16434 37214
rect 22878 37202 22930 37214
rect 30270 37202 30322 37214
rect 30718 37266 30770 37278
rect 30718 37202 30770 37214
rect 31166 37266 31218 37278
rect 31166 37202 31218 37214
rect 31390 37266 31442 37278
rect 31390 37202 31442 37214
rect 31726 37266 31778 37278
rect 31726 37202 31778 37214
rect 14030 37154 14082 37166
rect 13570 37102 13582 37154
rect 13634 37102 13646 37154
rect 14030 37090 14082 37102
rect 14814 37154 14866 37166
rect 16606 37154 16658 37166
rect 23662 37154 23714 37166
rect 15698 37102 15710 37154
rect 15762 37102 15774 37154
rect 19618 37102 19630 37154
rect 19682 37102 19694 37154
rect 14814 37090 14866 37102
rect 16606 37090 16658 37102
rect 23662 37090 23714 37102
rect 25566 37154 25618 37166
rect 25566 37090 25618 37102
rect 9550 37042 9602 37054
rect 9550 36978 9602 36990
rect 9886 37042 9938 37054
rect 9886 36978 9938 36990
rect 17278 37042 17330 37054
rect 17278 36978 17330 36990
rect 1344 36874 40544 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40544 36874
rect 1344 36788 40544 36822
rect 14926 36706 14978 36718
rect 27010 36654 27022 36706
rect 27074 36654 27086 36706
rect 14926 36642 14978 36654
rect 13806 36594 13858 36606
rect 8194 36542 8206 36594
rect 8258 36542 8270 36594
rect 10322 36542 10334 36594
rect 10386 36542 10398 36594
rect 12114 36542 12126 36594
rect 12178 36542 12190 36594
rect 13806 36530 13858 36542
rect 15150 36594 15202 36606
rect 15150 36530 15202 36542
rect 16942 36594 16994 36606
rect 16942 36530 16994 36542
rect 24894 36594 24946 36606
rect 26462 36594 26514 36606
rect 25778 36542 25790 36594
rect 25842 36542 25854 36594
rect 24894 36530 24946 36542
rect 26462 36530 26514 36542
rect 13582 36482 13634 36494
rect 7522 36430 7534 36482
rect 7586 36430 7598 36482
rect 12002 36430 12014 36482
rect 12066 36430 12078 36482
rect 13582 36418 13634 36430
rect 13694 36482 13746 36494
rect 13694 36418 13746 36430
rect 14030 36482 14082 36494
rect 14030 36418 14082 36430
rect 16046 36482 16098 36494
rect 16046 36418 16098 36430
rect 16718 36482 16770 36494
rect 16718 36418 16770 36430
rect 17838 36482 17890 36494
rect 20750 36482 20802 36494
rect 19394 36430 19406 36482
rect 19458 36430 19470 36482
rect 20178 36430 20190 36482
rect 20242 36430 20254 36482
rect 17838 36418 17890 36430
rect 20750 36418 20802 36430
rect 21534 36482 21586 36494
rect 21534 36418 21586 36430
rect 21646 36482 21698 36494
rect 21646 36418 21698 36430
rect 21758 36482 21810 36494
rect 21758 36418 21810 36430
rect 21870 36482 21922 36494
rect 26686 36482 26738 36494
rect 25442 36430 25454 36482
rect 25506 36430 25518 36482
rect 29362 36430 29374 36482
rect 29426 36430 29438 36482
rect 21870 36418 21922 36430
rect 26686 36418 26738 36430
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 12686 36370 12738 36382
rect 12686 36306 12738 36318
rect 15822 36370 15874 36382
rect 18946 36318 18958 36370
rect 19010 36318 19022 36370
rect 29138 36318 29150 36370
rect 29202 36318 29214 36370
rect 15822 36306 15874 36318
rect 12238 36258 12290 36270
rect 12238 36194 12290 36206
rect 12462 36258 12514 36270
rect 12462 36194 12514 36206
rect 13918 36258 13970 36270
rect 17166 36258 17218 36270
rect 14578 36206 14590 36258
rect 14642 36206 14654 36258
rect 16370 36206 16382 36258
rect 16434 36206 16446 36258
rect 13918 36194 13970 36206
rect 17166 36194 17218 36206
rect 17278 36258 17330 36270
rect 17278 36194 17330 36206
rect 17390 36258 17442 36270
rect 21422 36258 21474 36270
rect 18162 36206 18174 36258
rect 18226 36206 18238 36258
rect 17390 36194 17442 36206
rect 21422 36194 21474 36206
rect 22542 36258 22594 36270
rect 22542 36194 22594 36206
rect 31278 36258 31330 36270
rect 31278 36194 31330 36206
rect 1344 36090 40544 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40544 36090
rect 1344 36004 40544 36038
rect 15934 35922 15986 35934
rect 8418 35870 8430 35922
rect 8482 35870 8494 35922
rect 15934 35858 15986 35870
rect 17726 35922 17778 35934
rect 20850 35870 20862 35922
rect 20914 35870 20926 35922
rect 23314 35870 23326 35922
rect 23378 35870 23390 35922
rect 17726 35858 17778 35870
rect 9774 35810 9826 35822
rect 15710 35810 15762 35822
rect 9986 35758 9998 35810
rect 10050 35758 10062 35810
rect 11666 35758 11678 35810
rect 11730 35758 11742 35810
rect 9774 35746 9826 35758
rect 15710 35746 15762 35758
rect 16494 35810 16546 35822
rect 16494 35746 16546 35758
rect 16606 35810 16658 35822
rect 16606 35746 16658 35758
rect 17390 35810 17442 35822
rect 17390 35746 17442 35758
rect 17502 35810 17554 35822
rect 31502 35810 31554 35822
rect 30370 35758 30382 35810
rect 30434 35758 30446 35810
rect 32274 35758 32286 35810
rect 32338 35758 32350 35810
rect 17502 35746 17554 35758
rect 31502 35746 31554 35758
rect 13694 35698 13746 35710
rect 8194 35646 8206 35698
rect 8258 35646 8270 35698
rect 11218 35646 11230 35698
rect 11282 35646 11294 35698
rect 13694 35634 13746 35646
rect 15598 35698 15650 35710
rect 15598 35634 15650 35646
rect 20526 35698 20578 35710
rect 31278 35698 31330 35710
rect 33070 35698 33122 35710
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 26786 35646 26798 35698
rect 26850 35646 26862 35698
rect 32498 35646 32510 35698
rect 32562 35646 32574 35698
rect 20526 35634 20578 35646
rect 31278 35634 31330 35646
rect 33070 35634 33122 35646
rect 8878 35586 8930 35598
rect 8878 35522 8930 35534
rect 13470 35586 13522 35598
rect 13470 35522 13522 35534
rect 18062 35586 18114 35598
rect 18062 35522 18114 35534
rect 22990 35586 23042 35598
rect 22990 35522 23042 35534
rect 24782 35586 24834 35598
rect 33182 35586 33234 35598
rect 32162 35534 32174 35586
rect 32226 35534 32238 35586
rect 24782 35522 24834 35534
rect 33182 35522 33234 35534
rect 16494 35474 16546 35486
rect 14018 35422 14030 35474
rect 14082 35422 14094 35474
rect 16494 35410 16546 35422
rect 30942 35474 30994 35486
rect 30942 35410 30994 35422
rect 1344 35306 40544 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40544 35306
rect 1344 35220 40544 35254
rect 11678 35138 11730 35150
rect 11678 35074 11730 35086
rect 16830 35026 16882 35038
rect 27246 35026 27298 35038
rect 11218 34974 11230 35026
rect 11282 34974 11294 35026
rect 15250 34974 15262 35026
rect 15314 34974 15326 35026
rect 25890 34974 25902 35026
rect 25954 34974 25966 35026
rect 34514 34974 34526 35026
rect 34578 34974 34590 35026
rect 16830 34962 16882 34974
rect 27246 34962 27298 34974
rect 10782 34914 10834 34926
rect 19742 34914 19794 34926
rect 26238 34914 26290 34926
rect 10210 34862 10222 34914
rect 10274 34862 10286 34914
rect 12002 34862 12014 34914
rect 12066 34862 12078 34914
rect 14690 34862 14702 34914
rect 14754 34862 14766 34914
rect 23090 34862 23102 34914
rect 23154 34862 23166 34914
rect 26674 34862 26686 34914
rect 26738 34862 26750 34914
rect 30818 34862 30830 34914
rect 30882 34862 30894 34914
rect 31602 34862 31614 34914
rect 31666 34862 31678 34914
rect 10782 34850 10834 34862
rect 19742 34850 19794 34862
rect 26238 34850 26290 34862
rect 18846 34802 18898 34814
rect 10434 34750 10446 34802
rect 10498 34750 10510 34802
rect 18846 34738 18898 34750
rect 18958 34802 19010 34814
rect 18958 34738 19010 34750
rect 19406 34802 19458 34814
rect 30494 34802 30546 34814
rect 23762 34750 23774 34802
rect 23826 34750 23838 34802
rect 32386 34750 32398 34802
rect 32450 34750 32462 34802
rect 19406 34738 19458 34750
rect 30494 34738 30546 34750
rect 11790 34690 11842 34702
rect 11790 34626 11842 34638
rect 14926 34690 14978 34702
rect 14926 34626 14978 34638
rect 15150 34690 15202 34702
rect 15150 34626 15202 34638
rect 15262 34690 15314 34702
rect 15262 34626 15314 34638
rect 16382 34690 16434 34702
rect 16382 34626 16434 34638
rect 19182 34690 19234 34702
rect 19182 34626 19234 34638
rect 19518 34690 19570 34702
rect 19518 34626 19570 34638
rect 29934 34690 29986 34702
rect 29934 34626 29986 34638
rect 30158 34690 30210 34702
rect 30158 34626 30210 34638
rect 30382 34690 30434 34702
rect 30382 34626 30434 34638
rect 31054 34690 31106 34702
rect 31054 34626 31106 34638
rect 31278 34690 31330 34702
rect 31278 34626 31330 34638
rect 31390 34690 31442 34702
rect 31390 34626 31442 34638
rect 1344 34522 40544 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40544 34522
rect 1344 34436 40544 34470
rect 7870 34354 7922 34366
rect 7870 34290 7922 34302
rect 9774 34354 9826 34366
rect 9774 34290 9826 34302
rect 13246 34354 13298 34366
rect 16270 34354 16322 34366
rect 13570 34302 13582 34354
rect 13634 34302 13646 34354
rect 15698 34302 15710 34354
rect 15762 34302 15774 34354
rect 13246 34290 13298 34302
rect 16270 34290 16322 34302
rect 23438 34354 23490 34366
rect 23438 34290 23490 34302
rect 23886 34354 23938 34366
rect 23886 34290 23938 34302
rect 30494 34354 30546 34366
rect 30494 34290 30546 34302
rect 31278 34354 31330 34366
rect 31278 34290 31330 34302
rect 12014 34242 12066 34254
rect 8978 34190 8990 34242
rect 9042 34190 9054 34242
rect 12014 34178 12066 34190
rect 16046 34242 16098 34254
rect 16046 34178 16098 34190
rect 16494 34242 16546 34254
rect 30270 34242 30322 34254
rect 19506 34190 19518 34242
rect 19570 34190 19582 34242
rect 25778 34190 25790 34242
rect 25842 34190 25854 34242
rect 29698 34190 29710 34242
rect 29762 34190 29774 34242
rect 16494 34178 16546 34190
rect 30270 34178 30322 34190
rect 31054 34242 31106 34254
rect 31054 34178 31106 34190
rect 31390 34242 31442 34254
rect 31390 34178 31442 34190
rect 33070 34242 33122 34254
rect 33070 34178 33122 34190
rect 9662 34130 9714 34142
rect 8754 34078 8766 34130
rect 8818 34078 8830 34130
rect 9662 34066 9714 34078
rect 9886 34130 9938 34142
rect 9886 34066 9938 34078
rect 10334 34130 10386 34142
rect 10334 34066 10386 34078
rect 10558 34130 10610 34142
rect 10558 34066 10610 34078
rect 11790 34130 11842 34142
rect 11790 34066 11842 34078
rect 12126 34130 12178 34142
rect 12126 34066 12178 34078
rect 15374 34130 15426 34142
rect 15374 34066 15426 34078
rect 16606 34130 16658 34142
rect 16606 34066 16658 34078
rect 19182 34130 19234 34142
rect 19182 34066 19234 34078
rect 20190 34130 20242 34142
rect 20190 34066 20242 34078
rect 20302 34130 20354 34142
rect 20302 34066 20354 34078
rect 20526 34130 20578 34142
rect 20526 34066 20578 34078
rect 23662 34130 23714 34142
rect 23662 34066 23714 34078
rect 24110 34130 24162 34142
rect 24110 34066 24162 34078
rect 24334 34130 24386 34142
rect 24334 34066 24386 34078
rect 26126 34130 26178 34142
rect 26126 34066 26178 34078
rect 29038 34130 29090 34142
rect 29038 34066 29090 34078
rect 29374 34130 29426 34142
rect 29374 34066 29426 34078
rect 30158 34130 30210 34142
rect 30158 34066 30210 34078
rect 30942 34130 30994 34142
rect 30942 34066 30994 34078
rect 32286 34130 32338 34142
rect 33966 34130 34018 34142
rect 33506 34078 33518 34130
rect 33570 34078 33582 34130
rect 32286 34066 32338 34078
rect 33966 34066 34018 34078
rect 14254 34018 14306 34030
rect 10882 33966 10894 34018
rect 10946 33966 10958 34018
rect 14254 33954 14306 33966
rect 15150 34018 15202 34030
rect 15150 33954 15202 33966
rect 16382 34018 16434 34030
rect 16382 33954 16434 33966
rect 31838 34018 31890 34030
rect 31838 33954 31890 33966
rect 7758 33906 7810 33918
rect 7758 33842 7810 33854
rect 8094 33906 8146 33918
rect 8094 33842 8146 33854
rect 20638 33906 20690 33918
rect 31602 33854 31614 33906
rect 31666 33903 31678 33906
rect 31826 33903 31838 33906
rect 31666 33857 31838 33903
rect 31666 33854 31678 33857
rect 31826 33854 31838 33857
rect 31890 33854 31902 33906
rect 20638 33842 20690 33854
rect 1344 33738 40544 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40544 33738
rect 1344 33652 40544 33686
rect 13806 33570 13858 33582
rect 13806 33506 13858 33518
rect 18622 33570 18674 33582
rect 18622 33506 18674 33518
rect 32174 33570 32226 33582
rect 32174 33506 32226 33518
rect 11006 33458 11058 33470
rect 14926 33458 14978 33470
rect 5618 33406 5630 33458
rect 5682 33406 5694 33458
rect 7746 33406 7758 33458
rect 7810 33406 7822 33458
rect 9202 33406 9214 33458
rect 9266 33406 9278 33458
rect 13458 33406 13470 33458
rect 13522 33406 13534 33458
rect 11006 33394 11058 33406
rect 14926 33394 14978 33406
rect 15374 33458 15426 33470
rect 28478 33458 28530 33470
rect 15810 33406 15822 33458
rect 15874 33406 15886 33458
rect 20066 33406 20078 33458
rect 20130 33406 20142 33458
rect 27906 33406 27918 33458
rect 27970 33406 27982 33458
rect 30258 33406 30270 33458
rect 30322 33406 30334 33458
rect 15374 33394 15426 33406
rect 28478 33394 28530 33406
rect 11118 33346 11170 33358
rect 8530 33294 8542 33346
rect 8594 33294 8606 33346
rect 9538 33294 9550 33346
rect 9602 33294 9614 33346
rect 11118 33282 11170 33294
rect 11342 33346 11394 33358
rect 11342 33282 11394 33294
rect 14814 33346 14866 33358
rect 14814 33282 14866 33294
rect 15038 33346 15090 33358
rect 18398 33346 18450 33358
rect 16034 33294 16046 33346
rect 16098 33294 16110 33346
rect 15038 33282 15090 33294
rect 18398 33282 18450 33294
rect 19294 33346 19346 33358
rect 35198 33346 35250 33358
rect 19294 33282 19346 33294
rect 19630 33290 19682 33302
rect 25106 33294 25118 33346
rect 25170 33294 25182 33346
rect 30370 33294 30382 33346
rect 30434 33294 30446 33346
rect 8878 33234 8930 33246
rect 8878 33170 8930 33182
rect 10670 33234 10722 33246
rect 10670 33170 10722 33182
rect 11566 33234 11618 33246
rect 11566 33170 11618 33182
rect 11678 33234 11730 33246
rect 11678 33170 11730 33182
rect 13582 33234 13634 33246
rect 13582 33170 13634 33182
rect 14478 33234 14530 33246
rect 14478 33170 14530 33182
rect 19518 33234 19570 33246
rect 35198 33282 35250 33294
rect 19630 33226 19682 33238
rect 32286 33234 32338 33246
rect 19842 33182 19854 33234
rect 19906 33182 19918 33234
rect 22082 33182 22094 33234
rect 22146 33182 22158 33234
rect 25778 33182 25790 33234
rect 25842 33182 25854 33234
rect 29250 33182 29262 33234
rect 29314 33182 29326 33234
rect 19518 33170 19570 33182
rect 32286 33170 32338 33182
rect 34974 33234 35026 33246
rect 34974 33170 35026 33182
rect 35870 33234 35922 33246
rect 35870 33170 35922 33182
rect 36206 33234 36258 33246
rect 36206 33170 36258 33182
rect 10894 33122 10946 33134
rect 10894 33058 10946 33070
rect 16830 33122 16882 33134
rect 22430 33122 22482 33134
rect 18946 33070 18958 33122
rect 19010 33070 19022 33122
rect 16830 33058 16882 33070
rect 22430 33058 22482 33070
rect 31166 33122 31218 33134
rect 31166 33058 31218 33070
rect 31278 33122 31330 33134
rect 31278 33058 31330 33070
rect 31390 33122 31442 33134
rect 31390 33058 31442 33070
rect 31614 33122 31666 33134
rect 31614 33058 31666 33070
rect 32174 33122 32226 33134
rect 32174 33058 32226 33070
rect 35646 33122 35698 33134
rect 35646 33058 35698 33070
rect 35758 33122 35810 33134
rect 35758 33058 35810 33070
rect 36318 33122 36370 33134
rect 36318 33058 36370 33070
rect 36542 33122 36594 33134
rect 36542 33058 36594 33070
rect 37102 33122 37154 33134
rect 37102 33058 37154 33070
rect 1344 32954 40544 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40544 32954
rect 1344 32868 40544 32902
rect 8542 32786 8594 32798
rect 8542 32722 8594 32734
rect 8766 32786 8818 32798
rect 8766 32722 8818 32734
rect 23998 32786 24050 32798
rect 23998 32722 24050 32734
rect 25678 32786 25730 32798
rect 25678 32722 25730 32734
rect 26014 32786 26066 32798
rect 26014 32722 26066 32734
rect 26910 32786 26962 32798
rect 26910 32722 26962 32734
rect 27358 32786 27410 32798
rect 27358 32722 27410 32734
rect 29934 32786 29986 32798
rect 29934 32722 29986 32734
rect 33294 32786 33346 32798
rect 33294 32722 33346 32734
rect 37102 32786 37154 32798
rect 37102 32722 37154 32734
rect 8318 32674 8370 32686
rect 7634 32622 7646 32674
rect 7698 32622 7710 32674
rect 8318 32610 8370 32622
rect 10558 32674 10610 32686
rect 10558 32610 10610 32622
rect 17726 32674 17778 32686
rect 17726 32610 17778 32622
rect 19070 32674 19122 32686
rect 19070 32610 19122 32622
rect 19630 32674 19682 32686
rect 19630 32610 19682 32622
rect 24334 32674 24386 32686
rect 24334 32610 24386 32622
rect 24558 32674 24610 32686
rect 24558 32610 24610 32622
rect 28926 32674 28978 32686
rect 28926 32610 28978 32622
rect 29486 32674 29538 32686
rect 37774 32674 37826 32686
rect 31826 32622 31838 32674
rect 31890 32622 31902 32674
rect 33618 32622 33630 32674
rect 33682 32622 33694 32674
rect 29486 32610 29538 32622
rect 37774 32610 37826 32622
rect 7982 32562 8034 32574
rect 9662 32562 9714 32574
rect 17390 32562 17442 32574
rect 19406 32562 19458 32574
rect 8978 32510 8990 32562
rect 9042 32510 9054 32562
rect 10098 32510 10110 32562
rect 10162 32510 10174 32562
rect 16482 32510 16494 32562
rect 16546 32510 16558 32562
rect 18610 32510 18622 32562
rect 18674 32510 18686 32562
rect 18834 32510 18846 32562
rect 18898 32510 18910 32562
rect 7982 32498 8034 32510
rect 9662 32498 9714 32510
rect 17390 32498 17442 32510
rect 19406 32498 19458 32510
rect 19966 32562 20018 32574
rect 19966 32498 20018 32510
rect 20526 32562 20578 32574
rect 25566 32562 25618 32574
rect 20738 32510 20750 32562
rect 20802 32510 20814 32562
rect 20526 32498 20578 32510
rect 25566 32498 25618 32510
rect 25790 32562 25842 32574
rect 25790 32498 25842 32510
rect 29038 32562 29090 32574
rect 29038 32498 29090 32510
rect 29262 32562 29314 32574
rect 29262 32498 29314 32510
rect 29822 32562 29874 32574
rect 29822 32498 29874 32510
rect 30046 32562 30098 32574
rect 30046 32498 30098 32510
rect 30494 32562 30546 32574
rect 36878 32562 36930 32574
rect 37662 32562 37714 32574
rect 31042 32510 31054 32562
rect 31106 32510 31118 32562
rect 31378 32510 31390 32562
rect 31442 32510 31454 32562
rect 34402 32510 34414 32562
rect 34466 32510 34478 32562
rect 35970 32510 35982 32562
rect 36034 32510 36046 32562
rect 36642 32510 36654 32562
rect 36706 32510 36718 32562
rect 37314 32510 37326 32562
rect 37378 32510 37390 32562
rect 30494 32498 30546 32510
rect 36878 32498 36930 32510
rect 37662 32498 37714 32510
rect 8654 32450 8706 32462
rect 19854 32450 19906 32462
rect 33966 32450 34018 32462
rect 35310 32450 35362 32462
rect 36990 32450 37042 32462
rect 12226 32398 12238 32450
rect 12290 32398 12302 32450
rect 24658 32398 24670 32450
rect 24722 32398 24734 32450
rect 31490 32398 31502 32450
rect 31554 32398 31566 32450
rect 34738 32398 34750 32450
rect 34802 32398 34814 32450
rect 35634 32398 35646 32450
rect 35698 32398 35710 32450
rect 8654 32386 8706 32398
rect 19854 32386 19906 32398
rect 33966 32386 34018 32398
rect 35310 32386 35362 32398
rect 36990 32386 37042 32398
rect 19182 32338 19234 32350
rect 20626 32286 20638 32338
rect 20690 32286 20702 32338
rect 19182 32274 19234 32286
rect 1344 32170 40544 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40544 32170
rect 1344 32084 40544 32118
rect 12798 31890 12850 31902
rect 37886 31890 37938 31902
rect 15810 31838 15822 31890
rect 15874 31838 15886 31890
rect 18722 31838 18734 31890
rect 18786 31838 18798 31890
rect 34626 31838 34638 31890
rect 34690 31838 34702 31890
rect 12798 31826 12850 31838
rect 37886 31826 37938 31838
rect 16606 31778 16658 31790
rect 19742 31778 19794 31790
rect 15698 31726 15710 31778
rect 15762 31726 15774 31778
rect 18498 31726 18510 31778
rect 18562 31726 18574 31778
rect 16606 31714 16658 31726
rect 19742 31714 19794 31726
rect 23214 31778 23266 31790
rect 23214 31714 23266 31726
rect 23550 31778 23602 31790
rect 23550 31714 23602 31726
rect 24110 31778 24162 31790
rect 24110 31714 24162 31726
rect 24670 31778 24722 31790
rect 24670 31714 24722 31726
rect 26574 31778 26626 31790
rect 27582 31778 27634 31790
rect 33742 31778 33794 31790
rect 36206 31778 36258 31790
rect 27122 31726 27134 31778
rect 27186 31726 27198 31778
rect 28130 31726 28142 31778
rect 28194 31726 28206 31778
rect 31378 31726 31390 31778
rect 31442 31726 31454 31778
rect 33394 31726 33406 31778
rect 33458 31726 33470 31778
rect 34178 31726 34190 31778
rect 34242 31726 34254 31778
rect 35746 31726 35758 31778
rect 35810 31726 35822 31778
rect 26574 31714 26626 31726
rect 27582 31714 27634 31726
rect 33742 31714 33794 31726
rect 36206 31714 36258 31726
rect 36878 31778 36930 31790
rect 36878 31714 36930 31726
rect 37102 31778 37154 31790
rect 37102 31714 37154 31726
rect 37214 31778 37266 31790
rect 38210 31726 38222 31778
rect 38274 31726 38286 31778
rect 37214 31714 37266 31726
rect 12686 31666 12738 31678
rect 12686 31602 12738 31614
rect 19182 31666 19234 31678
rect 19182 31602 19234 31614
rect 20302 31666 20354 31678
rect 20302 31602 20354 31614
rect 21422 31666 21474 31678
rect 21422 31602 21474 31614
rect 21534 31666 21586 31678
rect 21534 31602 21586 31614
rect 23774 31666 23826 31678
rect 27470 31666 27522 31678
rect 25330 31614 25342 31666
rect 25394 31614 25406 31666
rect 23774 31602 23826 31614
rect 27470 31602 27522 31614
rect 30830 31666 30882 31678
rect 35310 31666 35362 31678
rect 33282 31614 33294 31666
rect 33346 31614 33358 31666
rect 30830 31602 30882 31614
rect 35310 31602 35362 31614
rect 37550 31666 37602 31678
rect 37550 31602 37602 31614
rect 8318 31554 8370 31566
rect 8318 31490 8370 31502
rect 9214 31554 9266 31566
rect 9214 31490 9266 31502
rect 20078 31554 20130 31566
rect 20078 31490 20130 31502
rect 20414 31554 20466 31566
rect 20414 31490 20466 31502
rect 20862 31554 20914 31566
rect 20862 31490 20914 31502
rect 21198 31554 21250 31566
rect 21198 31490 21250 31502
rect 21870 31554 21922 31566
rect 23550 31554 23602 31566
rect 22194 31502 22206 31554
rect 22258 31502 22270 31554
rect 21870 31490 21922 31502
rect 23550 31490 23602 31502
rect 25006 31554 25058 31566
rect 25006 31490 25058 31502
rect 25902 31554 25954 31566
rect 25902 31490 25954 31502
rect 26686 31554 26738 31566
rect 26686 31490 26738 31502
rect 26798 31554 26850 31566
rect 37998 31554 38050 31566
rect 29810 31502 29822 31554
rect 29874 31502 29886 31554
rect 26798 31490 26850 31502
rect 37998 31490 38050 31502
rect 38670 31554 38722 31566
rect 38670 31490 38722 31502
rect 1344 31386 40544 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40544 31386
rect 1344 31300 40544 31334
rect 19070 31218 19122 31230
rect 11666 31166 11678 31218
rect 11730 31166 11742 31218
rect 19070 31154 19122 31166
rect 26462 31218 26514 31230
rect 35534 31218 35586 31230
rect 26898 31166 26910 31218
rect 26962 31215 26974 31218
rect 27234 31215 27246 31218
rect 26962 31169 27246 31215
rect 26962 31166 26974 31169
rect 27234 31166 27246 31169
rect 27298 31166 27310 31218
rect 26462 31154 26514 31166
rect 35534 31154 35586 31166
rect 35870 31218 35922 31230
rect 35870 31154 35922 31166
rect 36542 31218 36594 31230
rect 36542 31154 36594 31166
rect 26238 31106 26290 31118
rect 12898 31054 12910 31106
rect 12962 31054 12974 31106
rect 25890 31054 25902 31106
rect 25954 31054 25966 31106
rect 26238 31042 26290 31054
rect 35086 31106 35138 31118
rect 35086 31042 35138 31054
rect 35310 31106 35362 31118
rect 37986 31054 37998 31106
rect 38050 31054 38062 31106
rect 35310 31042 35362 31054
rect 10110 30994 10162 31006
rect 15934 30994 15986 31006
rect 19182 30994 19234 31006
rect 24334 30994 24386 31006
rect 11442 30942 11454 30994
rect 11506 30942 11518 30994
rect 12226 30942 12238 30994
rect 12290 30942 12302 30994
rect 16370 30942 16382 30994
rect 16434 30942 16446 30994
rect 23874 30942 23886 30994
rect 23938 30942 23950 30994
rect 10110 30930 10162 30942
rect 15934 30930 15986 30942
rect 19182 30930 19234 30942
rect 24334 30930 24386 30942
rect 25566 30994 25618 31006
rect 25566 30930 25618 30942
rect 26798 30994 26850 31006
rect 35758 30994 35810 31006
rect 27234 30942 27246 30994
rect 27298 30942 27310 30994
rect 36306 30942 36318 30994
rect 36370 30942 36382 30994
rect 37202 30942 37214 30994
rect 37266 30942 37278 30994
rect 26798 30930 26850 30942
rect 35758 30930 35810 30942
rect 16830 30882 16882 30894
rect 15026 30830 15038 30882
rect 15090 30830 15102 30882
rect 16830 30818 16882 30830
rect 17502 30882 17554 30894
rect 35646 30882 35698 30894
rect 30258 30830 30270 30882
rect 30322 30830 30334 30882
rect 40114 30830 40126 30882
rect 40178 30830 40190 30882
rect 17502 30818 17554 30830
rect 35646 30818 35698 30830
rect 9886 30770 9938 30782
rect 9538 30718 9550 30770
rect 9602 30718 9614 30770
rect 9886 30706 9938 30718
rect 19070 30770 19122 30782
rect 19070 30706 19122 30718
rect 26574 30770 26626 30782
rect 26574 30706 26626 30718
rect 36654 30770 36706 30782
rect 36654 30706 36706 30718
rect 1344 30602 40544 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40544 30602
rect 1344 30516 40544 30550
rect 27582 30434 27634 30446
rect 27582 30370 27634 30382
rect 27806 30434 27858 30446
rect 27806 30370 27858 30382
rect 37662 30434 37714 30446
rect 37662 30370 37714 30382
rect 8206 30322 8258 30334
rect 8206 30258 8258 30270
rect 8990 30322 9042 30334
rect 8990 30258 9042 30270
rect 10894 30322 10946 30334
rect 30718 30322 30770 30334
rect 22978 30270 22990 30322
rect 23042 30270 23054 30322
rect 10894 30258 10946 30270
rect 30718 30258 30770 30270
rect 31278 30322 31330 30334
rect 32398 30322 32450 30334
rect 32050 30270 32062 30322
rect 32114 30270 32126 30322
rect 31278 30258 31330 30270
rect 32398 30258 32450 30270
rect 34638 30322 34690 30334
rect 34638 30258 34690 30270
rect 36318 30322 36370 30334
rect 37986 30270 37998 30322
rect 38050 30270 38062 30322
rect 36318 30258 36370 30270
rect 17838 30210 17890 30222
rect 8530 30158 8542 30210
rect 8594 30158 8606 30210
rect 9538 30158 9550 30210
rect 9602 30158 9614 30210
rect 9874 30158 9886 30210
rect 9938 30158 9950 30210
rect 17838 30146 17890 30158
rect 17950 30210 18002 30222
rect 17950 30146 18002 30158
rect 18174 30210 18226 30222
rect 18174 30146 18226 30158
rect 18398 30210 18450 30222
rect 23326 30210 23378 30222
rect 22754 30158 22766 30210
rect 22818 30158 22830 30210
rect 18398 30146 18450 30158
rect 23326 30146 23378 30158
rect 25902 30210 25954 30222
rect 25902 30146 25954 30158
rect 26462 30210 26514 30222
rect 26462 30146 26514 30158
rect 27134 30210 27186 30222
rect 27134 30146 27186 30158
rect 28030 30210 28082 30222
rect 28030 30146 28082 30158
rect 28366 30210 28418 30222
rect 31838 30210 31890 30222
rect 29250 30158 29262 30210
rect 29314 30158 29326 30210
rect 28366 30146 28418 30158
rect 31838 30146 31890 30158
rect 32958 30210 33010 30222
rect 32958 30146 33010 30158
rect 33966 30210 34018 30222
rect 33966 30146 34018 30158
rect 37326 30210 37378 30222
rect 37326 30146 37378 30158
rect 7870 30098 7922 30110
rect 18734 30098 18786 30110
rect 9986 30046 9998 30098
rect 10050 30046 10062 30098
rect 7870 30034 7922 30046
rect 18734 30034 18786 30046
rect 19182 30098 19234 30110
rect 19182 30034 19234 30046
rect 20862 30098 20914 30110
rect 26238 30098 26290 30110
rect 22194 30046 22206 30098
rect 22258 30046 22270 30098
rect 20862 30034 20914 30046
rect 26238 30034 26290 30046
rect 26910 30098 26962 30110
rect 30382 30098 30434 30110
rect 29474 30046 29486 30098
rect 29538 30046 29550 30098
rect 26910 30034 26962 30046
rect 30382 30034 30434 30046
rect 32174 30098 32226 30110
rect 32174 30034 32226 30046
rect 34414 30098 34466 30110
rect 34414 30034 34466 30046
rect 34526 30098 34578 30110
rect 36978 30046 36990 30098
rect 37042 30046 37054 30098
rect 34526 30034 34578 30046
rect 8094 29986 8146 29998
rect 8094 29922 8146 29934
rect 8318 29986 8370 29998
rect 12350 29986 12402 29998
rect 9426 29934 9438 29986
rect 9490 29934 9502 29986
rect 8318 29922 8370 29934
rect 12350 29922 12402 29934
rect 18510 29986 18562 29998
rect 18510 29922 18562 29934
rect 18622 29986 18674 29998
rect 18622 29922 18674 29934
rect 18958 29986 19010 29998
rect 18958 29922 19010 29934
rect 21534 29986 21586 29998
rect 21534 29922 21586 29934
rect 21870 29986 21922 29998
rect 21870 29922 21922 29934
rect 26014 29986 26066 29998
rect 26014 29922 26066 29934
rect 28478 29986 28530 29998
rect 28478 29922 28530 29934
rect 28702 29986 28754 29998
rect 28702 29922 28754 29934
rect 30606 29986 30658 29998
rect 30606 29922 30658 29934
rect 30830 29986 30882 29998
rect 30830 29922 30882 29934
rect 31166 29986 31218 29998
rect 31166 29922 31218 29934
rect 31390 29986 31442 29998
rect 31390 29922 31442 29934
rect 32622 29986 32674 29998
rect 32622 29922 32674 29934
rect 32846 29986 32898 29998
rect 35982 29986 36034 29998
rect 33618 29934 33630 29986
rect 33682 29934 33694 29986
rect 32846 29922 32898 29934
rect 35982 29922 36034 29934
rect 36430 29986 36482 29998
rect 36430 29922 36482 29934
rect 37886 29986 37938 29998
rect 37886 29922 37938 29934
rect 38446 29986 38498 29998
rect 38446 29922 38498 29934
rect 1344 29818 40544 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40544 29818
rect 1344 29732 40544 29766
rect 16718 29650 16770 29662
rect 16718 29586 16770 29598
rect 18958 29650 19010 29662
rect 18958 29586 19010 29598
rect 29598 29650 29650 29662
rect 29598 29586 29650 29598
rect 31950 29650 32002 29662
rect 31950 29586 32002 29598
rect 36094 29650 36146 29662
rect 36094 29586 36146 29598
rect 7982 29538 8034 29550
rect 7982 29474 8034 29486
rect 17502 29538 17554 29550
rect 21198 29538 21250 29550
rect 19282 29486 19294 29538
rect 19346 29486 19358 29538
rect 20738 29486 20750 29538
rect 20802 29486 20814 29538
rect 17502 29474 17554 29486
rect 21198 29474 21250 29486
rect 26574 29538 26626 29550
rect 26574 29474 26626 29486
rect 26910 29538 26962 29550
rect 26910 29474 26962 29486
rect 27022 29538 27074 29550
rect 27022 29474 27074 29486
rect 29486 29538 29538 29550
rect 31838 29538 31890 29550
rect 30594 29486 30606 29538
rect 30658 29486 30670 29538
rect 37986 29486 37998 29538
rect 38050 29486 38062 29538
rect 29486 29474 29538 29486
rect 31838 29474 31890 29486
rect 8878 29426 8930 29438
rect 8642 29374 8654 29426
rect 8706 29374 8718 29426
rect 8878 29362 8930 29374
rect 9662 29426 9714 29438
rect 9662 29362 9714 29374
rect 9774 29426 9826 29438
rect 9774 29362 9826 29374
rect 10222 29426 10274 29438
rect 16830 29426 16882 29438
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 10222 29362 10274 29374
rect 16830 29362 16882 29374
rect 17390 29426 17442 29438
rect 17390 29362 17442 29374
rect 18286 29426 18338 29438
rect 18286 29362 18338 29374
rect 18510 29426 18562 29438
rect 22766 29426 22818 29438
rect 19170 29374 19182 29426
rect 19234 29374 19246 29426
rect 20850 29374 20862 29426
rect 20914 29374 20926 29426
rect 21410 29374 21422 29426
rect 21474 29374 21486 29426
rect 21746 29374 21758 29426
rect 21810 29374 21822 29426
rect 18510 29362 18562 29374
rect 22766 29362 22818 29374
rect 23326 29426 23378 29438
rect 26686 29426 26738 29438
rect 33070 29426 33122 29438
rect 35534 29426 35586 29438
rect 24098 29374 24110 29426
rect 24162 29374 24174 29426
rect 30818 29374 30830 29426
rect 30882 29374 30894 29426
rect 33282 29374 33294 29426
rect 33346 29374 33358 29426
rect 35858 29374 35870 29426
rect 35922 29374 35934 29426
rect 37202 29374 37214 29426
rect 37266 29374 37278 29426
rect 23326 29362 23378 29374
rect 26686 29362 26738 29374
rect 33070 29362 33122 29374
rect 35534 29362 35586 29374
rect 9998 29314 10050 29326
rect 14478 29314 14530 29326
rect 10770 29262 10782 29314
rect 10834 29262 10846 29314
rect 12898 29262 12910 29314
rect 12962 29262 12974 29314
rect 9998 29250 10050 29262
rect 14478 29250 14530 29262
rect 18062 29314 18114 29326
rect 33854 29314 33906 29326
rect 36878 29314 36930 29326
rect 20066 29262 20078 29314
rect 20130 29262 20142 29314
rect 23762 29262 23774 29314
rect 23826 29262 23838 29314
rect 35970 29262 35982 29314
rect 36034 29262 36046 29314
rect 40114 29262 40126 29314
rect 40178 29262 40190 29314
rect 18062 29250 18114 29262
rect 33854 29250 33906 29262
rect 36878 29250 36930 29262
rect 16718 29202 16770 29214
rect 16718 29138 16770 29150
rect 17502 29202 17554 29214
rect 17502 29138 17554 29150
rect 29598 29202 29650 29214
rect 29598 29138 29650 29150
rect 1344 29034 40544 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40544 29034
rect 1344 28948 40544 28982
rect 5966 28866 6018 28878
rect 5966 28802 6018 28814
rect 19630 28866 19682 28878
rect 19630 28802 19682 28814
rect 19854 28866 19906 28878
rect 19854 28802 19906 28814
rect 9550 28754 9602 28766
rect 18062 28754 18114 28766
rect 5618 28702 5630 28754
rect 5682 28702 5694 28754
rect 7074 28702 7086 28754
rect 7138 28702 7150 28754
rect 9202 28702 9214 28754
rect 9266 28702 9278 28754
rect 10434 28702 10446 28754
rect 10498 28702 10510 28754
rect 11106 28702 11118 28754
rect 11170 28702 11182 28754
rect 15362 28702 15374 28754
rect 15426 28702 15438 28754
rect 17042 28702 17054 28754
rect 17106 28702 17118 28754
rect 9550 28690 9602 28702
rect 18062 28690 18114 28702
rect 24222 28754 24274 28766
rect 28478 28754 28530 28766
rect 25890 28702 25902 28754
rect 25954 28702 25966 28754
rect 28018 28702 28030 28754
rect 28082 28702 28094 28754
rect 31490 28702 31502 28754
rect 31554 28702 31566 28754
rect 24222 28690 24274 28702
rect 28478 28690 28530 28702
rect 13806 28642 13858 28654
rect 6290 28590 6302 28642
rect 6354 28590 6366 28642
rect 10210 28590 10222 28642
rect 10274 28590 10286 28642
rect 11554 28590 11566 28642
rect 11618 28590 11630 28642
rect 12562 28590 12574 28642
rect 12626 28590 12638 28642
rect 13806 28578 13858 28590
rect 13918 28642 13970 28654
rect 15710 28642 15762 28654
rect 18174 28642 18226 28654
rect 23662 28642 23714 28654
rect 14802 28590 14814 28642
rect 14866 28590 14878 28642
rect 16818 28590 16830 28642
rect 16882 28590 16894 28642
rect 18722 28590 18734 28642
rect 18786 28590 18798 28642
rect 19394 28590 19406 28642
rect 19458 28590 19470 28642
rect 13918 28578 13970 28590
rect 15710 28578 15762 28590
rect 18174 28578 18226 28590
rect 23662 28578 23714 28590
rect 24894 28642 24946 28654
rect 35422 28642 35474 28654
rect 25218 28590 25230 28642
rect 25282 28590 25294 28642
rect 31266 28590 31278 28642
rect 31330 28590 31342 28642
rect 24894 28578 24946 28590
rect 35422 28578 35474 28590
rect 38558 28642 38610 28654
rect 38558 28578 38610 28590
rect 12014 28530 12066 28542
rect 12014 28466 12066 28478
rect 13470 28530 13522 28542
rect 13470 28466 13522 28478
rect 14142 28530 14194 28542
rect 14142 28466 14194 28478
rect 14254 28530 14306 28542
rect 14254 28466 14306 28478
rect 17726 28530 17778 28542
rect 17726 28466 17778 28478
rect 31726 28530 31778 28542
rect 38210 28478 38222 28530
rect 38274 28478 38286 28530
rect 31726 28466 31778 28478
rect 5742 28418 5794 28430
rect 13582 28418 13634 28430
rect 12338 28366 12350 28418
rect 12402 28366 12414 28418
rect 5742 28354 5794 28366
rect 13582 28354 13634 28366
rect 19518 28418 19570 28430
rect 19518 28354 19570 28366
rect 22430 28418 22482 28430
rect 22430 28354 22482 28366
rect 24110 28418 24162 28430
rect 24110 28354 24162 28366
rect 24334 28418 24386 28430
rect 24334 28354 24386 28366
rect 35534 28418 35586 28430
rect 35534 28354 35586 28366
rect 35758 28418 35810 28430
rect 35758 28354 35810 28366
rect 1344 28250 40544 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40544 28250
rect 1344 28164 40544 28198
rect 9662 28082 9714 28094
rect 9662 28018 9714 28030
rect 18398 28082 18450 28094
rect 18398 28018 18450 28030
rect 33070 28082 33122 28094
rect 33070 28018 33122 28030
rect 17838 27970 17890 27982
rect 5394 27918 5406 27970
rect 5458 27918 5470 27970
rect 17838 27906 17890 27918
rect 18510 27970 18562 27982
rect 27358 27970 27410 27982
rect 32286 27970 32338 27982
rect 22530 27918 22542 27970
rect 22594 27918 22606 27970
rect 27906 27918 27918 27970
rect 27970 27918 27982 27970
rect 18510 27906 18562 27918
rect 27358 27906 27410 27918
rect 32286 27906 32338 27918
rect 9550 27858 9602 27870
rect 4722 27806 4734 27858
rect 4786 27806 4798 27858
rect 9550 27794 9602 27806
rect 9774 27858 9826 27870
rect 9774 27794 9826 27806
rect 10222 27858 10274 27870
rect 16382 27858 16434 27870
rect 18174 27858 18226 27870
rect 22878 27858 22930 27870
rect 28254 27858 28306 27870
rect 15922 27806 15934 27858
rect 15986 27806 15998 27858
rect 17490 27806 17502 27858
rect 17554 27806 17566 27858
rect 18834 27806 18846 27858
rect 18898 27806 18910 27858
rect 27570 27806 27582 27858
rect 27634 27806 27646 27858
rect 31826 27806 31838 27858
rect 31890 27806 31902 27858
rect 32050 27806 32062 27858
rect 32114 27806 32126 27858
rect 33282 27806 33294 27858
rect 33346 27806 33358 27858
rect 33506 27806 33518 27858
rect 33570 27806 33582 27858
rect 35858 27806 35870 27858
rect 35922 27806 35934 27858
rect 10222 27794 10274 27806
rect 16382 27794 16434 27806
rect 18174 27794 18226 27806
rect 22878 27794 22930 27806
rect 28254 27794 28306 27806
rect 19406 27746 19458 27758
rect 7522 27694 7534 27746
rect 7586 27694 7598 27746
rect 13346 27694 13358 27746
rect 13410 27694 13422 27746
rect 17602 27694 17614 27746
rect 17666 27694 17678 27746
rect 18946 27694 18958 27746
rect 19010 27694 19022 27746
rect 19406 27682 19458 27694
rect 25342 27746 25394 27758
rect 25342 27682 25394 27694
rect 35422 27746 35474 27758
rect 36306 27694 36318 27746
rect 36370 27694 36382 27746
rect 35422 27682 35474 27694
rect 27246 27634 27298 27646
rect 27246 27570 27298 27582
rect 31950 27634 32002 27646
rect 31950 27570 32002 27582
rect 32958 27634 33010 27646
rect 32958 27570 33010 27582
rect 1344 27466 40544 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40544 27466
rect 1344 27380 40544 27414
rect 17166 27298 17218 27310
rect 10322 27246 10334 27298
rect 10386 27295 10398 27298
rect 10994 27295 11006 27298
rect 10386 27249 11006 27295
rect 10386 27246 10398 27249
rect 10994 27246 11006 27249
rect 11058 27246 11070 27298
rect 17166 27234 17218 27246
rect 31950 27298 32002 27310
rect 31950 27234 32002 27246
rect 32174 27298 32226 27310
rect 32174 27234 32226 27246
rect 33854 27298 33906 27310
rect 35298 27246 35310 27298
rect 35362 27246 35374 27298
rect 37986 27246 37998 27298
rect 38050 27246 38062 27298
rect 33854 27234 33906 27246
rect 6974 27186 7026 27198
rect 6974 27122 7026 27134
rect 10558 27186 10610 27198
rect 10558 27122 10610 27134
rect 11006 27186 11058 27198
rect 12910 27186 12962 27198
rect 24670 27186 24722 27198
rect 26686 27186 26738 27198
rect 28030 27186 28082 27198
rect 12114 27134 12126 27186
rect 12178 27134 12190 27186
rect 15922 27134 15934 27186
rect 15986 27134 15998 27186
rect 18274 27134 18286 27186
rect 18338 27134 18350 27186
rect 21298 27134 21310 27186
rect 21362 27134 21374 27186
rect 25778 27134 25790 27186
rect 25842 27134 25854 27186
rect 27682 27134 27694 27186
rect 27746 27134 27758 27186
rect 11006 27122 11058 27134
rect 12910 27122 12962 27134
rect 24670 27122 24722 27134
rect 26686 27122 26738 27134
rect 28030 27122 28082 27134
rect 29822 27186 29874 27198
rect 32958 27186 33010 27198
rect 31602 27134 31614 27186
rect 31666 27134 31678 27186
rect 29822 27122 29874 27134
rect 32958 27122 33010 27134
rect 34862 27186 34914 27198
rect 38546 27134 38558 27186
rect 38610 27134 38622 27186
rect 34862 27122 34914 27134
rect 6526 27074 6578 27086
rect 16830 27074 16882 27086
rect 19294 27074 19346 27086
rect 12450 27022 12462 27074
rect 12514 27022 12526 27074
rect 16146 27022 16158 27074
rect 16210 27022 16222 27074
rect 17490 27022 17502 27074
rect 17554 27022 17566 27074
rect 6526 27010 6578 27022
rect 16830 27010 16882 27022
rect 19294 27010 19346 27022
rect 19518 27074 19570 27086
rect 19518 27010 19570 27022
rect 19742 27074 19794 27086
rect 20414 27074 20466 27086
rect 20178 27022 20190 27074
rect 20242 27022 20254 27074
rect 19742 27010 19794 27022
rect 20414 27010 20466 27022
rect 20638 27074 20690 27086
rect 29038 27074 29090 27086
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 26226 27022 26238 27074
rect 26290 27022 26302 27074
rect 27570 27022 27582 27074
rect 27634 27022 27646 27074
rect 20638 27010 20690 27022
rect 29038 27010 29090 27022
rect 29486 27074 29538 27086
rect 29486 27010 29538 27022
rect 29598 27074 29650 27086
rect 29598 27010 29650 27022
rect 30046 27074 30098 27086
rect 30046 27010 30098 27022
rect 31502 27074 31554 27086
rect 31502 27010 31554 27022
rect 32846 27074 32898 27086
rect 35422 27074 35474 27086
rect 39566 27074 39618 27086
rect 33282 27022 33294 27074
rect 33346 27022 33358 27074
rect 34290 27022 34302 27074
rect 34354 27022 34366 27074
rect 35970 27022 35982 27074
rect 36034 27022 36046 27074
rect 38322 27022 38334 27074
rect 38386 27022 38398 27074
rect 40002 27022 40014 27074
rect 40066 27022 40078 27074
rect 32846 27010 32898 27022
rect 35422 27010 35474 27022
rect 39566 27010 39618 27022
rect 18398 26962 18450 26974
rect 6178 26910 6190 26962
rect 6242 26910 6254 26962
rect 18398 26898 18450 26910
rect 18622 26962 18674 26974
rect 18622 26898 18674 26910
rect 20750 26962 20802 26974
rect 28590 26962 28642 26974
rect 23426 26910 23438 26962
rect 23490 26910 23502 26962
rect 20750 26898 20802 26910
rect 28590 26898 28642 26910
rect 31390 26962 31442 26974
rect 31390 26898 31442 26910
rect 33070 26962 33122 26974
rect 33070 26898 33122 26910
rect 34526 26962 34578 26974
rect 34738 26910 34750 26962
rect 34802 26910 34814 26962
rect 34526 26898 34578 26910
rect 17614 26850 17666 26862
rect 17614 26786 17666 26798
rect 17726 26850 17778 26862
rect 17726 26786 17778 26798
rect 17838 26850 17890 26862
rect 17838 26786 17890 26798
rect 19630 26850 19682 26862
rect 32734 26850 32786 26862
rect 29474 26798 29486 26850
rect 29538 26798 29550 26850
rect 19630 26786 19682 26798
rect 32734 26786 32786 26798
rect 39790 26850 39842 26862
rect 39790 26786 39842 26798
rect 1344 26682 40544 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40544 26682
rect 1344 26596 40544 26630
rect 19182 26514 19234 26526
rect 19182 26450 19234 26462
rect 19966 26514 20018 26526
rect 31390 26514 31442 26526
rect 39566 26514 39618 26526
rect 23538 26462 23550 26514
rect 23602 26462 23614 26514
rect 33282 26462 33294 26514
rect 33346 26462 33358 26514
rect 19966 26450 20018 26462
rect 31390 26450 31442 26462
rect 39566 26450 39618 26462
rect 3950 26402 4002 26414
rect 2034 26350 2046 26402
rect 2098 26350 2110 26402
rect 3950 26338 4002 26350
rect 19294 26402 19346 26414
rect 33070 26402 33122 26414
rect 28354 26350 28366 26402
rect 28418 26350 28430 26402
rect 19294 26338 19346 26350
rect 33070 26338 33122 26350
rect 34862 26402 34914 26414
rect 34862 26338 34914 26350
rect 36318 26402 36370 26414
rect 36318 26338 36370 26350
rect 39790 26402 39842 26414
rect 39790 26338 39842 26350
rect 40126 26402 40178 26414
rect 40126 26338 40178 26350
rect 23214 26290 23266 26302
rect 1810 26238 1822 26290
rect 1874 26238 1886 26290
rect 23214 26226 23266 26238
rect 24334 26290 24386 26302
rect 30942 26290 30994 26302
rect 27682 26238 27694 26290
rect 27746 26238 27758 26290
rect 24334 26226 24386 26238
rect 30942 26226 30994 26238
rect 31726 26290 31778 26302
rect 31726 26226 31778 26238
rect 32062 26290 32114 26302
rect 32062 26226 32114 26238
rect 32286 26290 32338 26302
rect 36430 26290 36482 26302
rect 33282 26238 33294 26290
rect 33346 26238 33358 26290
rect 33842 26238 33854 26290
rect 33906 26238 33918 26290
rect 35746 26238 35758 26290
rect 35810 26238 35822 26290
rect 36754 26238 36766 26290
rect 36818 26238 36830 26290
rect 32286 26226 32338 26238
rect 36430 26226 36482 26238
rect 2494 26178 2546 26190
rect 2494 26114 2546 26126
rect 20974 26178 21026 26190
rect 20974 26114 21026 26126
rect 24558 26178 24610 26190
rect 24558 26114 24610 26126
rect 26910 26178 26962 26190
rect 30482 26126 30494 26178
rect 30546 26126 30558 26178
rect 35298 26126 35310 26178
rect 35362 26126 35374 26178
rect 26910 26114 26962 26126
rect 3838 26066 3890 26078
rect 3838 26002 3890 26014
rect 4174 26066 4226 26078
rect 31502 26066 31554 26078
rect 23986 26014 23998 26066
rect 24050 26014 24062 26066
rect 30706 26014 30718 26066
rect 30770 26063 30782 26066
rect 31266 26063 31278 26066
rect 30770 26017 31278 26063
rect 30770 26014 30782 26017
rect 31266 26014 31278 26017
rect 31330 26014 31342 26066
rect 4174 26002 4226 26014
rect 31502 26002 31554 26014
rect 33518 26066 33570 26078
rect 33518 26002 33570 26014
rect 1344 25898 40544 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40544 25898
rect 1344 25812 40544 25846
rect 24334 25730 24386 25742
rect 24334 25666 24386 25678
rect 11454 25618 11506 25630
rect 23886 25618 23938 25630
rect 32958 25618 33010 25630
rect 34750 25618 34802 25630
rect 1698 25566 1710 25618
rect 1762 25566 1774 25618
rect 3826 25566 3838 25618
rect 3890 25566 3902 25618
rect 10322 25566 10334 25618
rect 10386 25566 10398 25618
rect 16370 25566 16382 25618
rect 16434 25566 16446 25618
rect 31154 25566 31166 25618
rect 31218 25566 31230 25618
rect 32162 25566 32174 25618
rect 32226 25566 32238 25618
rect 34066 25566 34078 25618
rect 34130 25566 34142 25618
rect 35634 25566 35646 25618
rect 35698 25566 35710 25618
rect 11454 25554 11506 25566
rect 23886 25554 23938 25566
rect 32958 25554 33010 25566
rect 34750 25554 34802 25566
rect 18846 25506 18898 25518
rect 30270 25506 30322 25518
rect 4610 25454 4622 25506
rect 4674 25454 4686 25506
rect 10098 25454 10110 25506
rect 10162 25454 10174 25506
rect 13458 25454 13470 25506
rect 13522 25454 13534 25506
rect 24770 25454 24782 25506
rect 24834 25454 24846 25506
rect 31042 25454 31054 25506
rect 31106 25454 31118 25506
rect 32498 25454 32510 25506
rect 32562 25454 32574 25506
rect 33730 25454 33742 25506
rect 33794 25454 33806 25506
rect 35186 25454 35198 25506
rect 35250 25454 35262 25506
rect 18846 25442 18898 25454
rect 30270 25442 30322 25454
rect 10894 25394 10946 25406
rect 22766 25394 22818 25406
rect 10210 25342 10222 25394
rect 10274 25342 10286 25394
rect 14242 25342 14254 25394
rect 14306 25342 14318 25394
rect 19170 25342 19182 25394
rect 19234 25342 19246 25394
rect 10894 25330 10946 25342
rect 22766 25330 22818 25342
rect 23774 25394 23826 25406
rect 23774 25330 23826 25342
rect 24222 25394 24274 25406
rect 31614 25394 31666 25406
rect 29474 25342 29486 25394
rect 29538 25391 29550 25394
rect 29698 25391 29710 25394
rect 29538 25345 29710 25391
rect 29538 25342 29550 25345
rect 29698 25342 29710 25345
rect 29762 25342 29774 25394
rect 29922 25342 29934 25394
rect 29986 25342 29998 25394
rect 24222 25330 24274 25342
rect 31614 25330 31666 25342
rect 33294 25394 33346 25406
rect 33294 25330 33346 25342
rect 9214 25282 9266 25294
rect 9214 25218 9266 25230
rect 11006 25282 11058 25294
rect 11006 25218 11058 25230
rect 22430 25282 22482 25294
rect 24994 25230 25006 25282
rect 25058 25230 25070 25282
rect 22430 25218 22482 25230
rect 1344 25114 40544 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40544 25114
rect 1344 25028 40544 25062
rect 6526 24946 6578 24958
rect 6526 24882 6578 24894
rect 10782 24946 10834 24958
rect 33406 24946 33458 24958
rect 31826 24894 31838 24946
rect 31890 24894 31902 24946
rect 10782 24882 10834 24894
rect 33406 24882 33458 24894
rect 33518 24946 33570 24958
rect 33518 24882 33570 24894
rect 33630 24946 33682 24958
rect 33630 24882 33682 24894
rect 36878 24946 36930 24958
rect 36878 24882 36930 24894
rect 6862 24834 6914 24846
rect 5282 24782 5294 24834
rect 5346 24782 5358 24834
rect 6862 24770 6914 24782
rect 22318 24834 22370 24846
rect 30818 24782 30830 24834
rect 30882 24782 30894 24834
rect 32274 24782 32286 24834
rect 32338 24782 32350 24834
rect 22318 24770 22370 24782
rect 6302 24722 6354 24734
rect 4610 24670 4622 24722
rect 4674 24670 4686 24722
rect 5058 24670 5070 24722
rect 5122 24670 5134 24722
rect 6302 24658 6354 24670
rect 6414 24722 6466 24734
rect 6414 24658 6466 24670
rect 6638 24722 6690 24734
rect 6638 24658 6690 24670
rect 7310 24722 7362 24734
rect 7310 24658 7362 24670
rect 7422 24722 7474 24734
rect 7422 24658 7474 24670
rect 7646 24722 7698 24734
rect 7646 24658 7698 24670
rect 7758 24722 7810 24734
rect 9774 24722 9826 24734
rect 8642 24670 8654 24722
rect 8706 24670 8718 24722
rect 7758 24658 7810 24670
rect 9774 24658 9826 24670
rect 10334 24722 10386 24734
rect 10334 24658 10386 24670
rect 10670 24722 10722 24734
rect 17502 24722 17554 24734
rect 11554 24670 11566 24722
rect 11618 24670 11630 24722
rect 10670 24658 10722 24670
rect 17502 24658 17554 24670
rect 17838 24722 17890 24734
rect 17838 24658 17890 24670
rect 18062 24722 18114 24734
rect 25790 24722 25842 24734
rect 21186 24670 21198 24722
rect 21250 24670 21262 24722
rect 22082 24670 22094 24722
rect 22146 24670 22158 24722
rect 18062 24658 18114 24670
rect 25790 24658 25842 24670
rect 26126 24722 26178 24734
rect 26126 24658 26178 24670
rect 26686 24722 26738 24734
rect 32958 24722 33010 24734
rect 31378 24670 31390 24722
rect 31442 24670 31454 24722
rect 32386 24670 32398 24722
rect 32450 24670 32462 24722
rect 37202 24670 37214 24722
rect 37266 24670 37278 24722
rect 26686 24658 26738 24670
rect 32958 24658 33010 24670
rect 7534 24610 7586 24622
rect 17614 24610 17666 24622
rect 25230 24610 25282 24622
rect 1698 24558 1710 24610
rect 1762 24558 1774 24610
rect 3826 24558 3838 24610
rect 3890 24558 3902 24610
rect 12338 24558 12350 24610
rect 12402 24558 12414 24610
rect 14466 24558 14478 24610
rect 14530 24558 14542 24610
rect 20850 24558 20862 24610
rect 20914 24558 20926 24610
rect 37986 24558 37998 24610
rect 38050 24558 38062 24610
rect 40114 24558 40126 24610
rect 40178 24558 40190 24610
rect 7534 24546 7586 24558
rect 17614 24546 17666 24558
rect 25230 24546 25282 24558
rect 8654 24498 8706 24510
rect 8654 24434 8706 24446
rect 8990 24498 9042 24510
rect 8990 24434 9042 24446
rect 10782 24498 10834 24510
rect 10782 24434 10834 24446
rect 1344 24330 40544 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40544 24330
rect 1344 24244 40544 24278
rect 3838 24162 3890 24174
rect 3838 24098 3890 24110
rect 4174 24162 4226 24174
rect 23874 24110 23886 24162
rect 23938 24110 23950 24162
rect 4174 24098 4226 24110
rect 18062 24050 18114 24062
rect 1922 23998 1934 24050
rect 1986 23998 1998 24050
rect 8530 23998 8542 24050
rect 8594 23998 8606 24050
rect 10658 23998 10670 24050
rect 10722 23998 10734 24050
rect 18062 23986 18114 23998
rect 18958 24050 19010 24062
rect 20750 24050 20802 24062
rect 20178 23998 20190 24050
rect 20242 23998 20254 24050
rect 40114 23998 40126 24050
rect 40178 23998 40190 24050
rect 18958 23986 19010 23998
rect 20750 23986 20802 23998
rect 6750 23938 6802 23950
rect 17054 23938 17106 23950
rect 2930 23886 2942 23938
rect 2994 23886 3006 23938
rect 3826 23886 3838 23938
rect 3890 23886 3902 23938
rect 7970 23886 7982 23938
rect 8034 23886 8046 23938
rect 11442 23886 11454 23938
rect 11506 23886 11518 23938
rect 16594 23886 16606 23938
rect 16658 23886 16670 23938
rect 6750 23874 6802 23886
rect 17054 23874 17106 23886
rect 17278 23938 17330 23950
rect 17278 23874 17330 23886
rect 17726 23938 17778 23950
rect 19854 23938 19906 23950
rect 23102 23938 23154 23950
rect 36542 23938 36594 23950
rect 18498 23886 18510 23938
rect 18562 23886 18574 23938
rect 22306 23886 22318 23938
rect 22370 23886 22382 23938
rect 23650 23886 23662 23938
rect 23714 23886 23726 23938
rect 24210 23886 24222 23938
rect 24274 23886 24286 23938
rect 37202 23886 37214 23938
rect 37266 23886 37278 23938
rect 17726 23874 17778 23886
rect 19854 23874 19906 23886
rect 23102 23874 23154 23886
rect 36542 23874 36594 23886
rect 6414 23826 6466 23838
rect 6414 23762 6466 23774
rect 19630 23826 19682 23838
rect 19630 23762 19682 23774
rect 20190 23826 20242 23838
rect 20190 23762 20242 23774
rect 20638 23826 20690 23838
rect 20638 23762 20690 23774
rect 22766 23826 22818 23838
rect 22766 23762 22818 23774
rect 24446 23826 24498 23838
rect 37986 23774 37998 23826
rect 38050 23774 38062 23826
rect 24446 23762 24498 23774
rect 6526 23714 6578 23726
rect 17502 23714 17554 23726
rect 7746 23662 7758 23714
rect 7810 23662 7822 23714
rect 16370 23662 16382 23714
rect 16434 23662 16446 23714
rect 6526 23650 6578 23662
rect 17502 23650 17554 23662
rect 17950 23714 18002 23726
rect 17950 23650 18002 23662
rect 18174 23714 18226 23726
rect 18174 23650 18226 23662
rect 20078 23714 20130 23726
rect 20078 23650 20130 23662
rect 21870 23714 21922 23726
rect 22878 23714 22930 23726
rect 22082 23662 22094 23714
rect 22146 23662 22158 23714
rect 21870 23650 21922 23662
rect 22878 23650 22930 23662
rect 24334 23714 24386 23726
rect 24334 23650 24386 23662
rect 29822 23714 29874 23726
rect 29822 23650 29874 23662
rect 1344 23546 40544 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40544 23546
rect 1344 23460 40544 23494
rect 4734 23378 4786 23390
rect 4734 23314 4786 23326
rect 5294 23378 5346 23390
rect 5294 23314 5346 23326
rect 6526 23378 6578 23390
rect 6526 23314 6578 23326
rect 7198 23378 7250 23390
rect 7198 23314 7250 23326
rect 36654 23378 36706 23390
rect 36654 23314 36706 23326
rect 37550 23378 37602 23390
rect 37550 23314 37602 23326
rect 4510 23266 4562 23278
rect 4510 23202 4562 23214
rect 5070 23266 5122 23278
rect 5070 23202 5122 23214
rect 5966 23266 6018 23278
rect 5966 23202 6018 23214
rect 7422 23266 7474 23278
rect 7422 23202 7474 23214
rect 8878 23266 8930 23278
rect 16382 23266 16434 23278
rect 15474 23214 15486 23266
rect 15538 23214 15550 23266
rect 8878 23202 8930 23214
rect 16382 23202 16434 23214
rect 18062 23266 18114 23278
rect 30046 23266 30098 23278
rect 23314 23214 23326 23266
rect 23378 23214 23390 23266
rect 18062 23202 18114 23214
rect 30046 23202 30098 23214
rect 34414 23266 34466 23278
rect 37438 23266 37490 23278
rect 36306 23214 36318 23266
rect 36370 23214 36382 23266
rect 34414 23202 34466 23214
rect 37438 23202 37490 23214
rect 4398 23154 4450 23166
rect 4398 23090 4450 23102
rect 4958 23154 5010 23166
rect 4958 23090 5010 23102
rect 5518 23154 5570 23166
rect 5518 23090 5570 23102
rect 5630 23154 5682 23166
rect 5630 23090 5682 23102
rect 5742 23154 5794 23166
rect 5742 23090 5794 23102
rect 7086 23154 7138 23166
rect 15822 23154 15874 23166
rect 10322 23102 10334 23154
rect 10386 23102 10398 23154
rect 12338 23102 12350 23154
rect 12402 23102 12414 23154
rect 13010 23102 13022 23154
rect 13074 23102 13086 23154
rect 7086 23090 7138 23102
rect 15822 23090 15874 23102
rect 16270 23154 16322 23166
rect 16270 23090 16322 23102
rect 17726 23154 17778 23166
rect 17726 23090 17778 23102
rect 17950 23154 18002 23166
rect 17950 23090 18002 23102
rect 18510 23154 18562 23166
rect 29822 23154 29874 23166
rect 19506 23102 19518 23154
rect 19570 23102 19582 23154
rect 26562 23102 26574 23154
rect 26626 23102 26638 23154
rect 18510 23090 18562 23102
rect 29822 23090 29874 23102
rect 30494 23154 30546 23166
rect 30494 23090 30546 23102
rect 34302 23154 34354 23166
rect 34302 23090 34354 23102
rect 34638 23154 34690 23166
rect 34638 23090 34690 23102
rect 9886 23042 9938 23054
rect 16158 23042 16210 23054
rect 15138 22990 15150 23042
rect 15202 22990 15214 23042
rect 9886 22978 9938 22990
rect 16158 22978 16210 22990
rect 19070 23042 19122 23054
rect 29934 23042 29986 23054
rect 27346 22990 27358 23042
rect 27410 22990 27422 23042
rect 29474 22990 29486 23042
rect 29538 22990 29550 23042
rect 19070 22978 19122 22990
rect 29934 22978 29986 22990
rect 6414 22930 6466 22942
rect 6414 22866 6466 22878
rect 6750 22930 6802 22942
rect 6750 22866 6802 22878
rect 8654 22930 8706 22942
rect 8654 22866 8706 22878
rect 8990 22930 9042 22942
rect 8990 22866 9042 22878
rect 17614 22930 17666 22942
rect 37662 22930 37714 22942
rect 18498 22878 18510 22930
rect 18562 22927 18574 22930
rect 18946 22927 18958 22930
rect 18562 22881 18958 22927
rect 18562 22878 18574 22881
rect 18946 22878 18958 22881
rect 19010 22878 19022 22930
rect 17614 22866 17666 22878
rect 37662 22866 37714 22878
rect 1344 22762 40544 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40544 22762
rect 1344 22676 40544 22710
rect 16494 22594 16546 22606
rect 16494 22530 16546 22542
rect 29038 22594 29090 22606
rect 29038 22530 29090 22542
rect 33742 22594 33794 22606
rect 33742 22530 33794 22542
rect 12126 22482 12178 22494
rect 28142 22482 28194 22494
rect 5058 22430 5070 22482
rect 5122 22430 5134 22482
rect 6402 22430 6414 22482
rect 6466 22430 6478 22482
rect 11330 22430 11342 22482
rect 11394 22430 11406 22482
rect 15698 22430 15710 22482
rect 15762 22430 15774 22482
rect 22978 22430 22990 22482
rect 23042 22430 23054 22482
rect 25106 22430 25118 22482
rect 25170 22430 25182 22482
rect 27346 22430 27358 22482
rect 27410 22430 27422 22482
rect 33394 22430 33406 22482
rect 33458 22430 33470 22482
rect 12126 22418 12178 22430
rect 28142 22418 28194 22430
rect 4734 22370 4786 22382
rect 15934 22370 15986 22382
rect 6290 22318 6302 22370
rect 6354 22318 6366 22370
rect 11666 22318 11678 22370
rect 11730 22318 11742 22370
rect 15362 22318 15374 22370
rect 15426 22318 15438 22370
rect 4734 22306 4786 22318
rect 15934 22306 15986 22318
rect 16270 22370 16322 22382
rect 16270 22306 16322 22318
rect 16718 22370 16770 22382
rect 16718 22306 16770 22318
rect 19630 22370 19682 22382
rect 19630 22306 19682 22318
rect 21646 22370 21698 22382
rect 26350 22370 26402 22382
rect 27806 22370 27858 22382
rect 37886 22370 37938 22382
rect 25778 22318 25790 22370
rect 25842 22318 25854 22370
rect 26786 22318 26798 22370
rect 26850 22318 26862 22370
rect 27458 22318 27470 22370
rect 27522 22318 27534 22370
rect 28242 22318 28254 22370
rect 28306 22318 28318 22370
rect 29362 22318 29374 22370
rect 29426 22318 29438 22370
rect 35298 22318 35310 22370
rect 35362 22318 35374 22370
rect 35858 22318 35870 22370
rect 35922 22318 35934 22370
rect 37314 22318 37326 22370
rect 37378 22318 37390 22370
rect 21646 22306 21698 22318
rect 26350 22306 26402 22318
rect 27806 22306 27858 22318
rect 37886 22306 37938 22318
rect 38222 22370 38274 22382
rect 38222 22306 38274 22318
rect 4958 22258 5010 22270
rect 28030 22258 28082 22270
rect 6178 22206 6190 22258
rect 6242 22206 6254 22258
rect 18274 22206 18286 22258
rect 18338 22206 18350 22258
rect 21298 22206 21310 22258
rect 21362 22206 21374 22258
rect 4958 22194 5010 22206
rect 28030 22194 28082 22206
rect 28478 22258 28530 22270
rect 28478 22194 28530 22206
rect 29598 22258 29650 22270
rect 29598 22194 29650 22206
rect 32734 22258 32786 22270
rect 32734 22194 32786 22206
rect 33070 22258 33122 22270
rect 33070 22194 33122 22206
rect 34190 22258 34242 22270
rect 34190 22194 34242 22206
rect 34414 22258 34466 22270
rect 36206 22258 36258 22270
rect 35522 22206 35534 22258
rect 35586 22206 35598 22258
rect 34414 22194 34466 22206
rect 36206 22194 36258 22206
rect 37998 22258 38050 22270
rect 37998 22194 38050 22206
rect 38558 22258 38610 22270
rect 38558 22194 38610 22206
rect 6526 22146 6578 22158
rect 6526 22082 6578 22094
rect 6750 22146 6802 22158
rect 6750 22082 6802 22094
rect 17166 22146 17218 22158
rect 17166 22082 17218 22094
rect 17950 22146 18002 22158
rect 27246 22146 27298 22158
rect 19282 22094 19294 22146
rect 19346 22094 19358 22146
rect 17950 22082 18002 22094
rect 27246 22082 27298 22094
rect 29150 22146 29202 22158
rect 29150 22082 29202 22094
rect 33518 22146 33570 22158
rect 33518 22082 33570 22094
rect 34526 22146 34578 22158
rect 34526 22082 34578 22094
rect 34638 22146 34690 22158
rect 34638 22082 34690 22094
rect 36094 22146 36146 22158
rect 36094 22082 36146 22094
rect 38446 22146 38498 22158
rect 38446 22082 38498 22094
rect 1344 21978 40544 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40544 21978
rect 1344 21892 40544 21926
rect 3054 21810 3106 21822
rect 3054 21746 3106 21758
rect 3502 21810 3554 21822
rect 5406 21810 5458 21822
rect 4834 21758 4846 21810
rect 4898 21758 4910 21810
rect 3502 21746 3554 21758
rect 5406 21746 5458 21758
rect 6750 21810 6802 21822
rect 6750 21746 6802 21758
rect 6862 21810 6914 21822
rect 6862 21746 6914 21758
rect 7198 21810 7250 21822
rect 7198 21746 7250 21758
rect 26910 21810 26962 21822
rect 26910 21746 26962 21758
rect 28926 21810 28978 21822
rect 36418 21758 36430 21810
rect 36482 21758 36494 21810
rect 37874 21758 37886 21810
rect 37938 21758 37950 21810
rect 28926 21746 28978 21758
rect 2942 21698 2994 21710
rect 6638 21698 6690 21710
rect 15374 21698 15426 21710
rect 3826 21646 3838 21698
rect 3890 21646 3902 21698
rect 7522 21646 7534 21698
rect 7586 21646 7598 21698
rect 13906 21646 13918 21698
rect 13970 21646 13982 21698
rect 2942 21634 2994 21646
rect 6638 21634 6690 21646
rect 15374 21634 15426 21646
rect 15710 21698 15762 21710
rect 15710 21634 15762 21646
rect 16382 21698 16434 21710
rect 16382 21634 16434 21646
rect 19294 21698 19346 21710
rect 19294 21634 19346 21646
rect 27918 21698 27970 21710
rect 27918 21634 27970 21646
rect 28142 21698 28194 21710
rect 28142 21634 28194 21646
rect 29598 21698 29650 21710
rect 29598 21634 29650 21646
rect 32174 21698 32226 21710
rect 32174 21634 32226 21646
rect 33070 21698 33122 21710
rect 33070 21634 33122 21646
rect 33406 21698 33458 21710
rect 37550 21698 37602 21710
rect 34850 21646 34862 21698
rect 34914 21646 34926 21698
rect 35186 21646 35198 21698
rect 35250 21646 35262 21698
rect 33406 21634 33458 21646
rect 37550 21634 37602 21646
rect 5182 21586 5234 21598
rect 6190 21586 6242 21598
rect 4610 21534 4622 21586
rect 4674 21534 4686 21586
rect 5618 21534 5630 21586
rect 5682 21534 5694 21586
rect 5954 21534 5966 21586
rect 6018 21534 6030 21586
rect 5182 21522 5234 21534
rect 6190 21522 6242 21534
rect 13582 21586 13634 21598
rect 13582 21522 13634 21534
rect 15262 21586 15314 21598
rect 15262 21522 15314 21534
rect 16158 21586 16210 21598
rect 16158 21522 16210 21534
rect 16270 21586 16322 21598
rect 16270 21522 16322 21534
rect 18174 21586 18226 21598
rect 27582 21586 27634 21598
rect 23762 21534 23774 21586
rect 23826 21534 23838 21586
rect 18174 21522 18226 21534
rect 27582 21522 27634 21534
rect 28814 21586 28866 21598
rect 28814 21522 28866 21534
rect 29486 21586 29538 21598
rect 32510 21586 32562 21598
rect 31490 21534 31502 21586
rect 31554 21534 31566 21586
rect 29486 21522 29538 21534
rect 32510 21522 32562 21534
rect 33182 21586 33234 21598
rect 33182 21522 33234 21534
rect 33630 21586 33682 21598
rect 35870 21586 35922 21598
rect 37214 21586 37266 21598
rect 35410 21534 35422 21586
rect 35474 21534 35486 21586
rect 36978 21534 36990 21586
rect 37042 21534 37054 21586
rect 38098 21534 38110 21586
rect 38162 21534 38174 21586
rect 39106 21534 39118 21586
rect 39170 21534 39182 21586
rect 33630 21522 33682 21534
rect 35870 21522 35922 21534
rect 37214 21522 37266 21534
rect 15598 21474 15650 21486
rect 17950 21474 18002 21486
rect 24222 21474 24274 21486
rect 5506 21422 5518 21474
rect 5570 21422 5582 21474
rect 16818 21422 16830 21474
rect 16882 21422 16894 21474
rect 19394 21422 19406 21474
rect 19458 21422 19470 21474
rect 20850 21422 20862 21474
rect 20914 21422 20926 21474
rect 22978 21422 22990 21474
rect 23042 21422 23054 21474
rect 15598 21410 15650 21422
rect 17950 21410 18002 21422
rect 24222 21410 24274 21422
rect 26126 21474 26178 21486
rect 26126 21410 26178 21422
rect 27694 21474 27746 21486
rect 27694 21410 27746 21422
rect 30158 21474 30210 21486
rect 30158 21410 30210 21422
rect 34190 21474 34242 21486
rect 40002 21422 40014 21474
rect 40066 21422 40078 21474
rect 34190 21410 34242 21422
rect 3054 21362 3106 21374
rect 3054 21298 3106 21310
rect 18398 21362 18450 21374
rect 18398 21298 18450 21310
rect 18846 21362 18898 21374
rect 18846 21298 18898 21310
rect 19070 21362 19122 21374
rect 19070 21298 19122 21310
rect 29598 21362 29650 21374
rect 29598 21298 29650 21310
rect 31502 21362 31554 21374
rect 31502 21298 31554 21310
rect 31838 21362 31890 21374
rect 31838 21298 31890 21310
rect 33854 21362 33906 21374
rect 33854 21298 33906 21310
rect 36094 21362 36146 21374
rect 36094 21298 36146 21310
rect 37438 21362 37490 21374
rect 37438 21298 37490 21310
rect 1344 21194 40544 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40544 21194
rect 1344 21108 40544 21142
rect 4958 21026 5010 21038
rect 4958 20962 5010 20974
rect 5742 21026 5794 21038
rect 5742 20962 5794 20974
rect 5854 21026 5906 21038
rect 21534 21026 21586 21038
rect 16706 20974 16718 21026
rect 16770 20974 16782 21026
rect 5854 20962 5906 20974
rect 21534 20962 21586 20974
rect 21870 21026 21922 21038
rect 21870 20962 21922 20974
rect 30830 21026 30882 21038
rect 30830 20962 30882 20974
rect 6862 20914 6914 20926
rect 12014 20914 12066 20926
rect 11666 20862 11678 20914
rect 11730 20862 11742 20914
rect 6862 20850 6914 20862
rect 12014 20850 12066 20862
rect 18846 20914 18898 20926
rect 40114 20862 40126 20914
rect 40178 20862 40190 20914
rect 18846 20850 18898 20862
rect 6078 20802 6130 20814
rect 3602 20750 3614 20802
rect 3666 20750 3678 20802
rect 6078 20738 6130 20750
rect 6190 20802 6242 20814
rect 12238 20802 12290 20814
rect 6626 20750 6638 20802
rect 6690 20750 6702 20802
rect 10098 20750 10110 20802
rect 10162 20750 10174 20802
rect 6190 20738 6242 20750
rect 12238 20738 12290 20750
rect 17278 20802 17330 20814
rect 18062 20802 18114 20814
rect 21758 20802 21810 20814
rect 17826 20750 17838 20802
rect 17890 20750 17902 20802
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 21298 20750 21310 20802
rect 21362 20750 21374 20802
rect 17278 20738 17330 20750
rect 18062 20738 18114 20750
rect 21758 20738 21810 20750
rect 29486 20802 29538 20814
rect 29486 20738 29538 20750
rect 29710 20802 29762 20814
rect 31502 20802 31554 20814
rect 31266 20750 31278 20802
rect 31330 20750 31342 20802
rect 29710 20738 29762 20750
rect 31502 20738 31554 20750
rect 31614 20802 31666 20814
rect 31614 20738 31666 20750
rect 31726 20802 31778 20814
rect 32162 20750 32174 20802
rect 32226 20750 32238 20802
rect 34178 20750 34190 20802
rect 34242 20750 34254 20802
rect 37202 20750 37214 20802
rect 37266 20750 37278 20802
rect 31726 20738 31778 20750
rect 1710 20690 1762 20702
rect 1710 20626 1762 20638
rect 3166 20690 3218 20702
rect 3166 20626 3218 20638
rect 5070 20690 5122 20702
rect 5070 20626 5122 20638
rect 6974 20690 7026 20702
rect 6974 20626 7026 20638
rect 9214 20690 9266 20702
rect 9214 20626 9266 20638
rect 9550 20690 9602 20702
rect 9550 20626 9602 20638
rect 11342 20690 11394 20702
rect 11342 20626 11394 20638
rect 11566 20690 11618 20702
rect 11566 20626 11618 20638
rect 13470 20690 13522 20702
rect 13470 20626 13522 20638
rect 13582 20690 13634 20702
rect 13582 20626 13634 20638
rect 16046 20690 16098 20702
rect 16046 20626 16098 20638
rect 16382 20690 16434 20702
rect 16382 20626 16434 20638
rect 17166 20690 17218 20702
rect 17166 20626 17218 20638
rect 17390 20690 17442 20702
rect 17390 20626 17442 20638
rect 18174 20690 18226 20702
rect 29150 20690 29202 20702
rect 19506 20638 19518 20690
rect 19570 20638 19582 20690
rect 19730 20638 19742 20690
rect 19794 20638 19806 20690
rect 18174 20626 18226 20638
rect 29150 20626 29202 20638
rect 33294 20690 33346 20702
rect 33294 20626 33346 20638
rect 34750 20690 34802 20702
rect 37986 20638 37998 20690
rect 38050 20638 38062 20690
rect 34750 20626 34802 20638
rect 2046 20578 2098 20590
rect 2046 20514 2098 20526
rect 2494 20578 2546 20590
rect 2494 20514 2546 20526
rect 2942 20578 2994 20590
rect 2942 20514 2994 20526
rect 3054 20578 3106 20590
rect 4174 20578 4226 20590
rect 4958 20578 5010 20590
rect 13806 20578 13858 20590
rect 29262 20578 29314 20590
rect 36430 20578 36482 20590
rect 3826 20526 3838 20578
rect 3890 20526 3902 20578
rect 4498 20526 4510 20578
rect 4562 20526 4574 20578
rect 9874 20526 9886 20578
rect 9938 20526 9950 20578
rect 12562 20526 12574 20578
rect 12626 20526 12638 20578
rect 18610 20526 18622 20578
rect 18674 20526 18686 20578
rect 33618 20526 33630 20578
rect 33682 20526 33694 20578
rect 3054 20514 3106 20526
rect 4174 20514 4226 20526
rect 4958 20514 5010 20526
rect 13806 20514 13858 20526
rect 29262 20514 29314 20526
rect 36430 20514 36482 20526
rect 1344 20410 40544 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40544 20410
rect 1344 20324 40544 20358
rect 5630 20242 5682 20254
rect 2370 20190 2382 20242
rect 2434 20190 2446 20242
rect 3826 20190 3838 20242
rect 3890 20190 3902 20242
rect 5630 20178 5682 20190
rect 5742 20242 5794 20254
rect 5742 20178 5794 20190
rect 6862 20242 6914 20254
rect 6862 20178 6914 20190
rect 8430 20242 8482 20254
rect 8430 20178 8482 20190
rect 17950 20242 18002 20254
rect 17950 20178 18002 20190
rect 18174 20242 18226 20254
rect 18174 20178 18226 20190
rect 20974 20242 21026 20254
rect 20974 20178 21026 20190
rect 25790 20242 25842 20254
rect 25790 20178 25842 20190
rect 33406 20242 33458 20254
rect 33406 20178 33458 20190
rect 34750 20242 34802 20254
rect 34750 20178 34802 20190
rect 6638 20130 6690 20142
rect 3266 20078 3278 20130
rect 3330 20078 3342 20130
rect 3714 20078 3726 20130
rect 3778 20078 3790 20130
rect 5282 20078 5294 20130
rect 5346 20078 5358 20130
rect 6638 20066 6690 20078
rect 11790 20130 11842 20142
rect 11790 20066 11842 20078
rect 12014 20130 12066 20142
rect 12014 20066 12066 20078
rect 13134 20130 13186 20142
rect 13134 20066 13186 20078
rect 13358 20130 13410 20142
rect 13358 20066 13410 20078
rect 13918 20130 13970 20142
rect 13918 20066 13970 20078
rect 14478 20130 14530 20142
rect 14478 20066 14530 20078
rect 14590 20130 14642 20142
rect 21646 20130 21698 20142
rect 19282 20078 19294 20130
rect 19346 20078 19358 20130
rect 20402 20078 20414 20130
rect 20466 20078 20478 20130
rect 14590 20066 14642 20078
rect 21646 20066 21698 20078
rect 26126 20130 26178 20142
rect 26126 20066 26178 20078
rect 27582 20130 27634 20142
rect 27582 20066 27634 20078
rect 34302 20130 34354 20142
rect 38894 20130 38946 20142
rect 34302 20066 34354 20078
rect 34638 20074 34690 20086
rect 4734 20018 4786 20030
rect 2146 19966 2158 20018
rect 2210 19966 2222 20018
rect 2706 19966 2718 20018
rect 2770 19966 2782 20018
rect 4274 19966 4286 20018
rect 4338 19966 4350 20018
rect 4734 19954 4786 19966
rect 5854 20018 5906 20030
rect 6526 20018 6578 20030
rect 6178 19966 6190 20018
rect 6242 19966 6254 20018
rect 5854 19954 5906 19966
rect 6526 19954 6578 19966
rect 8206 20018 8258 20030
rect 8206 19954 8258 19966
rect 8542 20018 8594 20030
rect 8542 19954 8594 19966
rect 8654 20018 8706 20030
rect 12798 20018 12850 20030
rect 8978 19966 8990 20018
rect 9042 19966 9054 20018
rect 10322 19966 10334 20018
rect 10386 19966 10398 20018
rect 12226 19966 12238 20018
rect 12290 19966 12302 20018
rect 12562 19966 12574 20018
rect 12626 19966 12638 20018
rect 8654 19954 8706 19966
rect 12798 19954 12850 19966
rect 13470 20018 13522 20030
rect 13470 19954 13522 19966
rect 13694 20018 13746 20030
rect 13694 19954 13746 19966
rect 14254 20018 14306 20030
rect 14254 19954 14306 19966
rect 17838 20018 17890 20030
rect 17838 19954 17890 19966
rect 19630 20018 19682 20030
rect 19630 19954 19682 19966
rect 20190 20018 20242 20030
rect 20190 19954 20242 19966
rect 20638 20018 20690 20030
rect 21198 20018 21250 20030
rect 20738 19966 20750 20018
rect 20802 19966 20814 20018
rect 20638 19954 20690 19966
rect 21198 19954 21250 19966
rect 21870 20018 21922 20030
rect 26686 20018 26738 20030
rect 29934 20018 29986 20030
rect 26338 19966 26350 20018
rect 26402 19966 26414 20018
rect 27234 19966 27246 20018
rect 27298 19966 27310 20018
rect 21870 19954 21922 19966
rect 26686 19954 26738 19966
rect 29934 19954 29986 19966
rect 31838 20018 31890 20030
rect 31838 19954 31890 19966
rect 32062 20018 32114 20030
rect 32062 19954 32114 19966
rect 32510 20018 32562 20030
rect 32510 19954 32562 19966
rect 33518 20018 33570 20030
rect 33518 19954 33570 19966
rect 33742 20018 33794 20030
rect 33742 19954 33794 19966
rect 34078 20018 34130 20030
rect 38894 20066 38946 20078
rect 39678 20130 39730 20142
rect 39678 20066 39730 20078
rect 34638 20010 34690 20022
rect 35086 20018 35138 20030
rect 34850 19966 34862 20018
rect 34914 19966 34926 20018
rect 35410 19966 35422 20018
rect 35474 19966 35486 20018
rect 37090 19966 37102 20018
rect 37154 19966 37166 20018
rect 34078 19954 34130 19966
rect 35086 19954 35138 19966
rect 9662 19906 9714 19918
rect 11006 19906 11058 19918
rect 18958 19906 19010 19918
rect 10098 19854 10110 19906
rect 10162 19854 10174 19906
rect 12002 19854 12014 19906
rect 12066 19854 12078 19906
rect 9662 19842 9714 19854
rect 11006 19842 11058 19854
rect 18958 19842 19010 19854
rect 21422 19906 21474 19918
rect 21422 19842 21474 19854
rect 25230 19906 25282 19918
rect 25230 19842 25282 19854
rect 26462 19906 26514 19918
rect 26462 19842 26514 19854
rect 27470 19906 27522 19918
rect 31266 19854 31278 19906
rect 31330 19854 31342 19906
rect 37314 19854 37326 19906
rect 37378 19854 37390 19906
rect 27470 19842 27522 19854
rect 14030 19794 14082 19806
rect 14030 19730 14082 19742
rect 32286 19794 32338 19806
rect 37874 19742 37886 19794
rect 37938 19742 37950 19794
rect 32286 19730 32338 19742
rect 1344 19626 40544 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40544 19626
rect 1344 19540 40544 19574
rect 3278 19458 3330 19470
rect 3278 19394 3330 19406
rect 5742 19458 5794 19470
rect 5742 19394 5794 19406
rect 10782 19458 10834 19470
rect 12014 19458 12066 19470
rect 11106 19406 11118 19458
rect 11170 19406 11182 19458
rect 10782 19394 10834 19406
rect 12014 19394 12066 19406
rect 12798 19458 12850 19470
rect 12798 19394 12850 19406
rect 15038 19458 15090 19470
rect 21422 19458 21474 19470
rect 20738 19406 20750 19458
rect 20802 19406 20814 19458
rect 15038 19394 15090 19406
rect 21422 19394 21474 19406
rect 23774 19458 23826 19470
rect 23774 19394 23826 19406
rect 37774 19458 37826 19470
rect 37774 19394 37826 19406
rect 2494 19346 2546 19358
rect 2494 19282 2546 19294
rect 3054 19346 3106 19358
rect 3054 19282 3106 19294
rect 4734 19346 4786 19358
rect 4734 19282 4786 19294
rect 9550 19346 9602 19358
rect 9550 19282 9602 19294
rect 10558 19346 10610 19358
rect 14478 19346 14530 19358
rect 13570 19294 13582 19346
rect 13634 19294 13646 19346
rect 21746 19294 21758 19346
rect 21810 19294 21822 19346
rect 28130 19294 28142 19346
rect 28194 19294 28206 19346
rect 37986 19294 37998 19346
rect 38050 19294 38062 19346
rect 40002 19294 40014 19346
rect 40066 19294 40078 19346
rect 10558 19282 10610 19294
rect 14478 19282 14530 19294
rect 1710 19234 1762 19246
rect 5630 19234 5682 19246
rect 4162 19182 4174 19234
rect 4226 19182 4238 19234
rect 4610 19182 4622 19234
rect 4674 19182 4686 19234
rect 1710 19170 1762 19182
rect 5630 19170 5682 19182
rect 7870 19234 7922 19246
rect 7870 19170 7922 19182
rect 8318 19234 8370 19246
rect 8318 19170 8370 19182
rect 8990 19234 9042 19246
rect 8990 19170 9042 19182
rect 9438 19234 9490 19246
rect 9438 19170 9490 19182
rect 12574 19234 12626 19246
rect 14814 19234 14866 19246
rect 18510 19234 18562 19246
rect 24334 19234 24386 19246
rect 14018 19182 14030 19234
rect 14082 19182 14094 19234
rect 15362 19182 15374 19234
rect 15426 19182 15438 19234
rect 18946 19182 18958 19234
rect 19010 19182 19022 19234
rect 19954 19182 19966 19234
rect 20018 19182 20030 19234
rect 12574 19170 12626 19182
rect 14814 19170 14866 19182
rect 18510 19170 18562 19182
rect 24334 19170 24386 19182
rect 24670 19234 24722 19246
rect 28590 19234 28642 19246
rect 32622 19234 32674 19246
rect 25218 19182 25230 19234
rect 25282 19182 25294 19234
rect 30370 19182 30382 19234
rect 30434 19182 30446 19234
rect 24670 19170 24722 19182
rect 28590 19170 28642 19182
rect 32622 19170 32674 19182
rect 37438 19234 37490 19246
rect 38882 19182 38894 19234
rect 38946 19182 38958 19234
rect 37438 19170 37490 19182
rect 2046 19122 2098 19134
rect 2046 19058 2098 19070
rect 6302 19122 6354 19134
rect 6302 19058 6354 19070
rect 7310 19122 7362 19134
rect 7310 19058 7362 19070
rect 7534 19122 7586 19134
rect 7534 19058 7586 19070
rect 9662 19122 9714 19134
rect 9662 19058 9714 19070
rect 12238 19122 12290 19134
rect 12238 19058 12290 19070
rect 17278 19122 17330 19134
rect 20190 19122 20242 19134
rect 17602 19070 17614 19122
rect 17666 19070 17678 19122
rect 18050 19070 18062 19122
rect 18114 19070 18126 19122
rect 19506 19070 19518 19122
rect 19570 19070 19582 19122
rect 17278 19058 17330 19070
rect 20190 19058 20242 19070
rect 20302 19122 20354 19134
rect 20302 19058 20354 19070
rect 21646 19122 21698 19134
rect 21646 19058 21698 19070
rect 23886 19122 23938 19134
rect 23886 19058 23938 19070
rect 24894 19122 24946 19134
rect 29486 19122 29538 19134
rect 26002 19070 26014 19122
rect 26066 19070 26078 19122
rect 24894 19058 24946 19070
rect 29486 19058 29538 19070
rect 30606 19122 30658 19134
rect 30606 19058 30658 19070
rect 31278 19122 31330 19134
rect 31278 19058 31330 19070
rect 31614 19122 31666 19134
rect 31614 19058 31666 19070
rect 32958 19122 33010 19134
rect 32958 19058 33010 19070
rect 6414 19010 6466 19022
rect 3602 18958 3614 19010
rect 3666 18958 3678 19010
rect 6414 18946 6466 18958
rect 6638 19010 6690 19022
rect 6638 18946 6690 18958
rect 7758 19010 7810 19022
rect 7758 18946 7810 18958
rect 8206 19010 8258 19022
rect 8206 18946 8258 18958
rect 8430 19010 8482 19022
rect 8430 18946 8482 18958
rect 8654 19010 8706 19022
rect 8654 18946 8706 18958
rect 12910 19010 12962 19022
rect 24782 19010 24834 19022
rect 19394 18958 19406 19010
rect 19458 18958 19470 19010
rect 12910 18946 12962 18958
rect 24782 18946 24834 18958
rect 29822 19010 29874 19022
rect 29822 18946 29874 18958
rect 30942 19010 30994 19022
rect 30942 18946 30994 18958
rect 31950 19010 32002 19022
rect 37998 19010 38050 19022
rect 37090 18958 37102 19010
rect 37154 18958 37166 19010
rect 31950 18946 32002 18958
rect 37998 18946 38050 18958
rect 1344 18842 40544 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40544 18842
rect 1344 18756 40544 18790
rect 3838 18674 3890 18686
rect 3838 18610 3890 18622
rect 4286 18674 4338 18686
rect 4286 18610 4338 18622
rect 5182 18674 5234 18686
rect 5182 18610 5234 18622
rect 5294 18674 5346 18686
rect 5294 18610 5346 18622
rect 7422 18674 7474 18686
rect 7422 18610 7474 18622
rect 8206 18674 8258 18686
rect 8206 18610 8258 18622
rect 8990 18674 9042 18686
rect 8990 18610 9042 18622
rect 13918 18674 13970 18686
rect 13918 18610 13970 18622
rect 18846 18674 18898 18686
rect 18846 18610 18898 18622
rect 20078 18674 20130 18686
rect 20078 18610 20130 18622
rect 20974 18674 21026 18686
rect 37326 18674 37378 18686
rect 33730 18622 33742 18674
rect 33794 18622 33806 18674
rect 20974 18610 21026 18622
rect 37326 18610 37378 18622
rect 6078 18562 6130 18574
rect 6078 18498 6130 18510
rect 6302 18562 6354 18574
rect 6302 18498 6354 18510
rect 7646 18562 7698 18574
rect 7646 18498 7698 18510
rect 12910 18562 12962 18574
rect 12910 18498 12962 18510
rect 13246 18562 13298 18574
rect 13246 18498 13298 18510
rect 14142 18562 14194 18574
rect 25566 18562 25618 18574
rect 19730 18510 19742 18562
rect 19794 18510 19806 18562
rect 14142 18498 14194 18510
rect 25566 18498 25618 18510
rect 26350 18562 26402 18574
rect 34638 18562 34690 18574
rect 29250 18510 29262 18562
rect 29314 18510 29326 18562
rect 26350 18498 26402 18510
rect 34638 18498 34690 18510
rect 36654 18562 36706 18574
rect 36654 18498 36706 18510
rect 3726 18450 3778 18462
rect 3726 18386 3778 18398
rect 4174 18450 4226 18462
rect 4174 18386 4226 18398
rect 4510 18450 4562 18462
rect 5854 18450 5906 18462
rect 7870 18450 7922 18462
rect 5506 18398 5518 18450
rect 5570 18398 5582 18450
rect 7186 18398 7198 18450
rect 7250 18398 7262 18450
rect 4510 18386 4562 18398
rect 5854 18386 5906 18398
rect 7870 18386 7922 18398
rect 8206 18450 8258 18462
rect 8206 18386 8258 18398
rect 8430 18450 8482 18462
rect 17838 18450 17890 18462
rect 13682 18398 13694 18450
rect 13746 18398 13758 18450
rect 8430 18386 8482 18398
rect 17838 18386 17890 18398
rect 18286 18450 18338 18462
rect 25342 18450 25394 18462
rect 21522 18398 21534 18450
rect 21586 18398 21598 18450
rect 22194 18398 22206 18450
rect 22258 18398 22270 18450
rect 18286 18386 18338 18398
rect 25342 18386 25394 18398
rect 26574 18450 26626 18462
rect 34078 18450 34130 18462
rect 27234 18398 27246 18450
rect 27298 18398 27310 18450
rect 26574 18386 26626 18398
rect 34078 18386 34130 18398
rect 34414 18450 34466 18462
rect 34414 18386 34466 18398
rect 35086 18450 35138 18462
rect 36542 18450 36594 18462
rect 36082 18398 36094 18450
rect 36146 18398 36158 18450
rect 35086 18386 35138 18398
rect 36542 18386 36594 18398
rect 38894 18450 38946 18462
rect 38894 18386 38946 18398
rect 39678 18450 39730 18462
rect 39678 18386 39730 18398
rect 7310 18338 7362 18350
rect 34862 18338 34914 18350
rect 24322 18286 24334 18338
rect 24386 18286 24398 18338
rect 25666 18286 25678 18338
rect 25730 18286 25742 18338
rect 7310 18274 7362 18286
rect 34862 18274 34914 18286
rect 35310 18338 35362 18350
rect 36318 18338 36370 18350
rect 35522 18286 35534 18338
rect 35586 18286 35598 18338
rect 35310 18274 35362 18286
rect 36318 18274 36370 18286
rect 6414 18226 6466 18238
rect 6414 18162 6466 18174
rect 14254 18226 14306 18238
rect 26910 18226 26962 18238
rect 18386 18174 18398 18226
rect 18450 18223 18462 18226
rect 18834 18223 18846 18226
rect 18450 18177 18846 18223
rect 18450 18174 18462 18177
rect 18834 18174 18846 18177
rect 18898 18174 18910 18226
rect 14254 18162 14306 18174
rect 26910 18162 26962 18174
rect 38110 18226 38162 18238
rect 38110 18162 38162 18174
rect 1344 18058 40544 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40544 18058
rect 1344 17972 40544 18006
rect 19070 17890 19122 17902
rect 17154 17838 17166 17890
rect 17218 17838 17230 17890
rect 17826 17838 17838 17890
rect 17890 17838 17902 17890
rect 34514 17838 34526 17890
rect 34578 17838 34590 17890
rect 19070 17826 19122 17838
rect 24558 17778 24610 17790
rect 19506 17726 19518 17778
rect 19570 17726 19582 17778
rect 24558 17714 24610 17726
rect 25006 17778 25058 17790
rect 25006 17714 25058 17726
rect 27022 17778 27074 17790
rect 27022 17714 27074 17726
rect 27470 17778 27522 17790
rect 35522 17726 35534 17778
rect 35586 17726 35598 17778
rect 37762 17726 37774 17778
rect 37826 17726 37838 17778
rect 27470 17714 27522 17726
rect 6862 17666 6914 17678
rect 5954 17614 5966 17666
rect 6018 17614 6030 17666
rect 6862 17602 6914 17614
rect 7198 17666 7250 17678
rect 18398 17666 18450 17678
rect 20078 17666 20130 17678
rect 16818 17614 16830 17666
rect 16882 17614 16894 17666
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 18610 17614 18622 17666
rect 18674 17614 18686 17666
rect 19730 17614 19742 17666
rect 19794 17614 19806 17666
rect 7198 17602 7250 17614
rect 18398 17602 18450 17614
rect 20078 17602 20130 17614
rect 27694 17666 27746 17678
rect 27694 17602 27746 17614
rect 28254 17666 28306 17678
rect 28254 17602 28306 17614
rect 29150 17666 29202 17678
rect 31838 17666 31890 17678
rect 30706 17614 30718 17666
rect 30770 17614 30782 17666
rect 29150 17602 29202 17614
rect 31838 17602 31890 17614
rect 32398 17666 32450 17678
rect 32398 17602 32450 17614
rect 33966 17666 34018 17678
rect 35634 17614 35646 17666
rect 35698 17614 35710 17666
rect 37090 17614 37102 17666
rect 37154 17614 37166 17666
rect 33966 17602 34018 17614
rect 6190 17554 6242 17566
rect 6190 17490 6242 17502
rect 6974 17554 7026 17566
rect 6974 17490 7026 17502
rect 16606 17554 16658 17566
rect 16606 17490 16658 17502
rect 18286 17554 18338 17566
rect 18286 17490 18338 17502
rect 18958 17554 19010 17566
rect 18958 17490 19010 17502
rect 19518 17554 19570 17566
rect 19518 17490 19570 17502
rect 27134 17554 27186 17566
rect 30158 17554 30210 17566
rect 27906 17502 27918 17554
rect 27970 17502 27982 17554
rect 27134 17490 27186 17502
rect 30158 17490 30210 17502
rect 30494 17554 30546 17566
rect 30494 17490 30546 17502
rect 31166 17554 31218 17566
rect 31166 17490 31218 17502
rect 31502 17554 31554 17566
rect 31502 17490 31554 17502
rect 32622 17554 32674 17566
rect 32622 17490 32674 17502
rect 32734 17554 32786 17566
rect 32734 17490 32786 17502
rect 33854 17554 33906 17566
rect 33854 17490 33906 17502
rect 34078 17554 34130 17566
rect 34078 17490 34130 17502
rect 36318 17554 36370 17566
rect 36318 17490 36370 17502
rect 16718 17442 16770 17454
rect 16718 17378 16770 17390
rect 26686 17442 26738 17454
rect 26686 17378 26738 17390
rect 28478 17442 28530 17454
rect 28478 17378 28530 17390
rect 29486 17442 29538 17454
rect 29486 17378 29538 17390
rect 29822 17442 29874 17454
rect 29822 17378 29874 17390
rect 32174 17442 32226 17454
rect 40002 17390 40014 17442
rect 40066 17390 40078 17442
rect 32174 17378 32226 17390
rect 1344 17274 40544 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40544 17274
rect 1344 17188 40544 17222
rect 4398 17106 4450 17118
rect 4398 17042 4450 17054
rect 6526 17106 6578 17118
rect 6526 17042 6578 17054
rect 16494 17106 16546 17118
rect 16494 17042 16546 17054
rect 33406 17106 33458 17118
rect 36766 17106 36818 17118
rect 34066 17054 34078 17106
rect 34130 17054 34142 17106
rect 33406 17042 33458 17054
rect 36766 17042 36818 17054
rect 5742 16994 5794 17006
rect 4722 16942 4734 16994
rect 4786 16942 4798 16994
rect 5742 16930 5794 16942
rect 6302 16994 6354 17006
rect 16718 16994 16770 17006
rect 15474 16942 15486 16994
rect 15538 16942 15550 16994
rect 6302 16930 6354 16942
rect 16718 16930 16770 16942
rect 17726 16994 17778 17006
rect 17726 16930 17778 16942
rect 29150 16994 29202 17006
rect 29150 16930 29202 16942
rect 29486 16994 29538 17006
rect 29486 16930 29538 16942
rect 30158 16994 30210 17006
rect 30158 16930 30210 16942
rect 30494 16994 30546 17006
rect 30494 16930 30546 16942
rect 30830 16994 30882 17006
rect 30830 16930 30882 16942
rect 33070 16994 33122 17006
rect 33070 16930 33122 16942
rect 36542 16994 36594 17006
rect 36542 16930 36594 16942
rect 36654 16994 36706 17006
rect 37986 16942 37998 16994
rect 38050 16942 38062 16994
rect 36654 16930 36706 16942
rect 5630 16882 5682 16894
rect 3266 16830 3278 16882
rect 3330 16830 3342 16882
rect 5630 16818 5682 16830
rect 5966 16882 6018 16894
rect 5966 16818 6018 16830
rect 6190 16882 6242 16894
rect 6190 16818 6242 16830
rect 7310 16882 7362 16894
rect 7310 16818 7362 16830
rect 7534 16882 7586 16894
rect 7534 16818 7586 16830
rect 7758 16882 7810 16894
rect 7758 16818 7810 16830
rect 8206 16882 8258 16894
rect 16830 16882 16882 16894
rect 34638 16882 34690 16894
rect 8754 16830 8766 16882
rect 8818 16830 8830 16882
rect 16258 16830 16270 16882
rect 16322 16830 16334 16882
rect 19618 16830 19630 16882
rect 19682 16830 19694 16882
rect 29922 16830 29934 16882
rect 29986 16830 29998 16882
rect 8206 16818 8258 16830
rect 16830 16818 16882 16830
rect 34638 16818 34690 16830
rect 34974 16882 35026 16894
rect 35522 16830 35534 16882
rect 35586 16830 35598 16882
rect 37202 16830 37214 16882
rect 37266 16830 37278 16882
rect 34974 16818 35026 16830
rect 7646 16770 7698 16782
rect 17950 16770 18002 16782
rect 34414 16770 34466 16782
rect 13346 16718 13358 16770
rect 13410 16718 13422 16770
rect 19282 16718 19294 16770
rect 19346 16718 19358 16770
rect 7646 16706 7698 16718
rect 17950 16706 18002 16718
rect 34414 16706 34466 16718
rect 35198 16770 35250 16782
rect 35198 16706 35250 16718
rect 36206 16770 36258 16782
rect 40114 16718 40126 16770
rect 40178 16718 40190 16770
rect 36206 16706 36258 16718
rect 3278 16658 3330 16670
rect 3278 16594 3330 16606
rect 3614 16658 3666 16670
rect 3614 16594 3666 16606
rect 7086 16658 7138 16670
rect 7086 16594 7138 16606
rect 8430 16658 8482 16670
rect 8430 16594 8482 16606
rect 18174 16658 18226 16670
rect 18174 16594 18226 16606
rect 18398 16658 18450 16670
rect 18398 16594 18450 16606
rect 18846 16658 18898 16670
rect 18846 16594 18898 16606
rect 1344 16490 40544 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40544 16490
rect 1344 16404 40544 16438
rect 5518 16322 5570 16334
rect 5518 16258 5570 16270
rect 6190 16322 6242 16334
rect 6190 16258 6242 16270
rect 6750 16322 6802 16334
rect 6750 16258 6802 16270
rect 7086 16322 7138 16334
rect 17950 16322 18002 16334
rect 16930 16270 16942 16322
rect 16994 16319 17006 16322
rect 17602 16319 17614 16322
rect 16994 16273 17614 16319
rect 16994 16270 17006 16273
rect 17602 16270 17614 16273
rect 17666 16270 17678 16322
rect 7086 16258 7138 16270
rect 17950 16258 18002 16270
rect 33518 16322 33570 16334
rect 33518 16258 33570 16270
rect 33854 16322 33906 16334
rect 33854 16258 33906 16270
rect 34638 16322 34690 16334
rect 34638 16258 34690 16270
rect 39678 16322 39730 16334
rect 39678 16258 39730 16270
rect 8542 16210 8594 16222
rect 2482 16158 2494 16210
rect 2546 16158 2558 16210
rect 4610 16158 4622 16210
rect 4674 16158 4686 16210
rect 7522 16158 7534 16210
rect 7586 16158 7598 16210
rect 8542 16146 8594 16158
rect 16494 16210 16546 16222
rect 16494 16146 16546 16158
rect 17054 16210 17106 16222
rect 17054 16146 17106 16158
rect 17614 16210 17666 16222
rect 22878 16210 22930 16222
rect 22418 16158 22430 16210
rect 22482 16158 22494 16210
rect 17614 16146 17666 16158
rect 22878 16146 22930 16158
rect 25566 16210 25618 16222
rect 38322 16158 38334 16210
rect 38386 16158 38398 16210
rect 25566 16146 25618 16158
rect 5966 16098 6018 16110
rect 1810 16046 1822 16098
rect 1874 16046 1886 16098
rect 5966 16034 6018 16046
rect 6414 16098 6466 16110
rect 6414 16034 6466 16046
rect 7870 16098 7922 16110
rect 9438 16098 9490 16110
rect 8082 16046 8094 16098
rect 8146 16046 8158 16098
rect 7870 16034 7922 16046
rect 9438 16034 9490 16046
rect 18958 16098 19010 16110
rect 18958 16034 19010 16046
rect 25118 16098 25170 16110
rect 25118 16034 25170 16046
rect 31614 16098 31666 16110
rect 31614 16034 31666 16046
rect 34302 16098 34354 16110
rect 34302 16034 34354 16046
rect 34526 16098 34578 16110
rect 38894 16098 38946 16110
rect 37314 16046 37326 16098
rect 37378 16046 37390 16098
rect 34526 16034 34578 16046
rect 38894 16034 38946 16046
rect 7646 15986 7698 15998
rect 7646 15922 7698 15934
rect 18286 15986 18338 15998
rect 18286 15922 18338 15934
rect 22094 15986 22146 15998
rect 22094 15922 22146 15934
rect 22318 15986 22370 15998
rect 22318 15922 22370 15934
rect 23438 15986 23490 15998
rect 23438 15922 23490 15934
rect 24334 15986 24386 15998
rect 24334 15922 24386 15934
rect 24670 15986 24722 15998
rect 24670 15922 24722 15934
rect 31950 15986 32002 15998
rect 31950 15922 32002 15934
rect 33742 15986 33794 15998
rect 33742 15922 33794 15934
rect 5070 15874 5122 15886
rect 5070 15810 5122 15822
rect 6974 15874 7026 15886
rect 6974 15810 7026 15822
rect 7534 15874 7586 15886
rect 18062 15874 18114 15886
rect 9762 15822 9774 15874
rect 9826 15822 9838 15874
rect 7534 15810 7586 15822
rect 18062 15810 18114 15822
rect 19294 15874 19346 15886
rect 19294 15810 19346 15822
rect 23326 15874 23378 15886
rect 23326 15810 23378 15822
rect 33182 15874 33234 15886
rect 33182 15810 33234 15822
rect 34638 15874 34690 15886
rect 34638 15810 34690 15822
rect 36430 15874 36482 15886
rect 36430 15810 36482 15822
rect 1344 15706 40544 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40544 15706
rect 1344 15620 40544 15654
rect 5630 15538 5682 15550
rect 5630 15474 5682 15486
rect 6190 15538 6242 15550
rect 6190 15474 6242 15486
rect 7758 15538 7810 15550
rect 7758 15474 7810 15486
rect 9774 15538 9826 15550
rect 9774 15474 9826 15486
rect 10782 15538 10834 15550
rect 10782 15474 10834 15486
rect 16382 15538 16434 15550
rect 16382 15474 16434 15486
rect 16830 15538 16882 15550
rect 16830 15474 16882 15486
rect 17950 15538 18002 15550
rect 17950 15474 18002 15486
rect 19742 15538 19794 15550
rect 19742 15474 19794 15486
rect 29822 15538 29874 15550
rect 29822 15474 29874 15486
rect 33406 15538 33458 15550
rect 33406 15474 33458 15486
rect 37326 15538 37378 15550
rect 37326 15474 37378 15486
rect 38894 15538 38946 15550
rect 38894 15474 38946 15486
rect 39678 15538 39730 15550
rect 39678 15474 39730 15486
rect 7646 15426 7698 15438
rect 7646 15362 7698 15374
rect 8430 15426 8482 15438
rect 8430 15362 8482 15374
rect 8990 15426 9042 15438
rect 14478 15426 14530 15438
rect 11890 15374 11902 15426
rect 11954 15374 11966 15426
rect 13682 15374 13694 15426
rect 13746 15374 13758 15426
rect 8990 15362 9042 15374
rect 14478 15362 14530 15374
rect 17726 15426 17778 15438
rect 17726 15362 17778 15374
rect 18174 15426 18226 15438
rect 29934 15426 29986 15438
rect 22530 15374 22542 15426
rect 22594 15374 22606 15426
rect 25666 15374 25678 15426
rect 25730 15374 25742 15426
rect 27234 15374 27246 15426
rect 27298 15374 27310 15426
rect 18174 15362 18226 15374
rect 29934 15362 29986 15374
rect 31614 15426 31666 15438
rect 31614 15362 31666 15374
rect 33070 15426 33122 15438
rect 33070 15362 33122 15374
rect 5518 15314 5570 15326
rect 5518 15250 5570 15262
rect 6078 15314 6130 15326
rect 6078 15250 6130 15262
rect 7198 15314 7250 15326
rect 7198 15250 7250 15262
rect 7870 15314 7922 15326
rect 7870 15250 7922 15262
rect 8766 15314 8818 15326
rect 8766 15250 8818 15262
rect 9662 15314 9714 15326
rect 9662 15250 9714 15262
rect 9886 15314 9938 15326
rect 9886 15250 9938 15262
rect 10334 15314 10386 15326
rect 10334 15250 10386 15262
rect 11566 15314 11618 15326
rect 19070 15314 19122 15326
rect 19630 15314 19682 15326
rect 13906 15262 13918 15314
rect 13970 15262 13982 15314
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 19394 15262 19406 15314
rect 19458 15262 19470 15314
rect 11566 15250 11618 15262
rect 19070 15250 19122 15262
rect 19630 15250 19682 15262
rect 19854 15314 19906 15326
rect 19854 15250 19906 15262
rect 19966 15314 20018 15326
rect 30494 15314 30546 15326
rect 21858 15262 21870 15314
rect 21922 15262 21934 15314
rect 30146 15262 30158 15314
rect 30210 15262 30222 15314
rect 19966 15250 20018 15262
rect 30494 15250 30546 15262
rect 30942 15314 30994 15326
rect 30942 15250 30994 15262
rect 31166 15314 31218 15326
rect 31166 15250 31218 15262
rect 31390 15314 31442 15326
rect 32162 15262 32174 15314
rect 32226 15262 32238 15314
rect 31390 15250 31442 15262
rect 8542 15202 8594 15214
rect 8542 15138 8594 15150
rect 15374 15202 15426 15214
rect 15374 15138 15426 15150
rect 18958 15202 19010 15214
rect 27470 15202 27522 15214
rect 24658 15150 24670 15202
rect 24722 15150 24734 15202
rect 25330 15150 25342 15202
rect 25394 15150 25406 15202
rect 38098 15150 38110 15202
rect 38162 15150 38174 15202
rect 18958 15138 19010 15150
rect 27470 15138 27522 15150
rect 5630 15090 5682 15102
rect 5630 15026 5682 15038
rect 6190 15090 6242 15102
rect 6190 15026 6242 15038
rect 14366 15090 14418 15102
rect 14366 15026 14418 15038
rect 18062 15090 18114 15102
rect 18062 15026 18114 15038
rect 18734 15090 18786 15102
rect 18734 15026 18786 15038
rect 31054 15090 31106 15102
rect 31054 15026 31106 15038
rect 32174 15090 32226 15102
rect 32174 15026 32226 15038
rect 32510 15090 32562 15102
rect 32510 15026 32562 15038
rect 1344 14922 40544 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40544 14922
rect 1344 14836 40544 14870
rect 16046 14754 16098 14766
rect 16046 14690 16098 14702
rect 16718 14754 16770 14766
rect 16718 14690 16770 14702
rect 18734 14754 18786 14766
rect 18734 14690 18786 14702
rect 4958 14642 5010 14654
rect 4958 14578 5010 14590
rect 5070 14642 5122 14654
rect 7086 14642 7138 14654
rect 21422 14642 21474 14654
rect 6178 14590 6190 14642
rect 6242 14590 6254 14642
rect 14578 14590 14590 14642
rect 14642 14590 14654 14642
rect 17826 14590 17838 14642
rect 17890 14590 17902 14642
rect 5070 14578 5122 14590
rect 7086 14578 7138 14590
rect 21422 14578 21474 14590
rect 23886 14642 23938 14654
rect 23886 14578 23938 14590
rect 29150 14642 29202 14654
rect 29150 14578 29202 14590
rect 30830 14642 30882 14654
rect 39554 14590 39566 14642
rect 39618 14590 39630 14642
rect 30830 14578 30882 14590
rect 6974 14530 7026 14542
rect 5954 14478 5966 14530
rect 6018 14478 6030 14530
rect 6974 14466 7026 14478
rect 12238 14530 12290 14542
rect 12238 14466 12290 14478
rect 12350 14530 12402 14542
rect 12350 14466 12402 14478
rect 12462 14530 12514 14542
rect 12910 14530 12962 14542
rect 15710 14530 15762 14542
rect 18958 14530 19010 14542
rect 12562 14478 12574 14530
rect 12626 14478 12638 14530
rect 14018 14478 14030 14530
rect 14082 14478 14094 14530
rect 14466 14478 14478 14530
rect 14530 14478 14542 14530
rect 18386 14478 18398 14530
rect 18450 14478 18462 14530
rect 12462 14466 12514 14478
rect 12910 14466 12962 14478
rect 15710 14466 15762 14478
rect 18958 14466 19010 14478
rect 19294 14530 19346 14542
rect 19294 14466 19346 14478
rect 20078 14530 20130 14542
rect 20078 14466 20130 14478
rect 20750 14530 20802 14542
rect 20750 14466 20802 14478
rect 22206 14530 22258 14542
rect 22206 14466 22258 14478
rect 22766 14530 22818 14542
rect 23774 14530 23826 14542
rect 23426 14478 23438 14530
rect 23490 14478 23502 14530
rect 22766 14466 22818 14478
rect 23774 14466 23826 14478
rect 23998 14530 24050 14542
rect 30046 14530 30098 14542
rect 38894 14530 38946 14542
rect 25106 14478 25118 14530
rect 25170 14478 25182 14530
rect 25890 14478 25902 14530
rect 25954 14478 25966 14530
rect 29810 14478 29822 14530
rect 29874 14478 29886 14530
rect 31154 14478 31166 14530
rect 31218 14478 31230 14530
rect 23998 14466 24050 14478
rect 30046 14466 30098 14478
rect 38894 14466 38946 14478
rect 4846 14418 4898 14430
rect 4846 14354 4898 14366
rect 6638 14418 6690 14430
rect 15374 14418 15426 14430
rect 13458 14366 13470 14418
rect 13522 14366 13534 14418
rect 15026 14366 15038 14418
rect 15090 14366 15102 14418
rect 6638 14354 6690 14366
rect 15374 14354 15426 14366
rect 16158 14418 16210 14430
rect 16158 14354 16210 14366
rect 16830 14418 16882 14430
rect 16830 14354 16882 14366
rect 17390 14418 17442 14430
rect 17390 14354 17442 14366
rect 17950 14418 18002 14430
rect 26574 14418 26626 14430
rect 19730 14366 19742 14418
rect 19794 14366 19806 14418
rect 24770 14366 24782 14418
rect 24834 14366 24846 14418
rect 36194 14366 36206 14418
rect 36258 14366 36270 14418
rect 17950 14354 18002 14366
rect 26574 14354 26626 14366
rect 15598 14306 15650 14318
rect 15598 14242 15650 14254
rect 16718 14306 16770 14318
rect 16718 14242 16770 14254
rect 17614 14306 17666 14318
rect 17614 14242 17666 14254
rect 17838 14306 17890 14318
rect 17838 14242 17890 14254
rect 18622 14306 18674 14318
rect 18622 14242 18674 14254
rect 19182 14306 19234 14318
rect 20402 14254 20414 14306
rect 20466 14254 20478 14306
rect 19182 14242 19234 14254
rect 1344 14138 40544 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40544 14138
rect 1344 14052 40544 14086
rect 5070 13970 5122 13982
rect 5070 13906 5122 13918
rect 6078 13970 6130 13982
rect 6078 13906 6130 13918
rect 8094 13970 8146 13982
rect 8094 13906 8146 13918
rect 8206 13970 8258 13982
rect 8206 13906 8258 13918
rect 8430 13970 8482 13982
rect 8430 13906 8482 13918
rect 9662 13970 9714 13982
rect 9662 13906 9714 13918
rect 13470 13970 13522 13982
rect 13470 13906 13522 13918
rect 15486 13970 15538 13982
rect 19406 13970 19458 13982
rect 18274 13918 18286 13970
rect 18338 13918 18350 13970
rect 15486 13906 15538 13918
rect 19406 13906 19458 13918
rect 20302 13970 20354 13982
rect 20302 13906 20354 13918
rect 20750 13970 20802 13982
rect 20750 13906 20802 13918
rect 25342 13970 25394 13982
rect 25342 13906 25394 13918
rect 25454 13970 25506 13982
rect 29822 13970 29874 13982
rect 28578 13918 28590 13970
rect 28642 13918 28654 13970
rect 25454 13906 25506 13918
rect 29822 13906 29874 13918
rect 30494 13970 30546 13982
rect 30494 13906 30546 13918
rect 30718 13970 30770 13982
rect 30718 13906 30770 13918
rect 5742 13858 5794 13870
rect 2482 13806 2494 13858
rect 2546 13806 2558 13858
rect 5742 13794 5794 13806
rect 5854 13858 5906 13870
rect 9998 13858 10050 13870
rect 16382 13858 16434 13870
rect 7522 13806 7534 13858
rect 7586 13855 7598 13858
rect 7858 13855 7870 13858
rect 7586 13809 7870 13855
rect 7586 13806 7598 13809
rect 7858 13806 7870 13809
rect 7922 13806 7934 13858
rect 11554 13806 11566 13858
rect 11618 13806 11630 13858
rect 12226 13806 12238 13858
rect 12290 13806 12302 13858
rect 5854 13794 5906 13806
rect 9998 13794 10050 13806
rect 16382 13794 16434 13806
rect 16830 13858 16882 13870
rect 19070 13858 19122 13870
rect 17938 13806 17950 13858
rect 18002 13806 18014 13858
rect 18162 13806 18174 13858
rect 18226 13806 18238 13858
rect 16830 13794 16882 13806
rect 19070 13794 19122 13806
rect 19182 13858 19234 13870
rect 19182 13794 19234 13806
rect 25678 13858 25730 13870
rect 30158 13858 30210 13870
rect 26898 13806 26910 13858
rect 26962 13806 26974 13858
rect 25678 13794 25730 13806
rect 30158 13794 30210 13806
rect 32174 13858 32226 13870
rect 35634 13806 35646 13858
rect 35698 13806 35710 13858
rect 32174 13794 32226 13806
rect 10334 13746 10386 13758
rect 15038 13746 15090 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 8642 13694 8654 13746
rect 8706 13694 8718 13746
rect 11442 13694 11454 13746
rect 11506 13694 11518 13746
rect 12002 13694 12014 13746
rect 12066 13694 12078 13746
rect 12898 13694 12910 13746
rect 12962 13694 12974 13746
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 10334 13682 10386 13694
rect 15038 13682 15090 13694
rect 15598 13746 15650 13758
rect 19854 13746 19906 13758
rect 15922 13694 15934 13746
rect 15986 13694 15998 13746
rect 16594 13694 16606 13746
rect 16658 13694 16670 13746
rect 17714 13694 17726 13746
rect 17778 13694 17790 13746
rect 15598 13682 15650 13694
rect 19854 13682 19906 13694
rect 25230 13746 25282 13758
rect 31166 13746 31218 13758
rect 27458 13694 27470 13746
rect 27522 13694 27534 13746
rect 28130 13694 28142 13746
rect 28194 13694 28206 13746
rect 25230 13682 25282 13694
rect 31166 13682 31218 13694
rect 31390 13746 31442 13758
rect 31390 13682 31442 13694
rect 31614 13746 31666 13758
rect 31614 13682 31666 13694
rect 32510 13746 32562 13758
rect 36418 13694 36430 13746
rect 36482 13694 36494 13746
rect 32510 13682 32562 13694
rect 8318 13634 8370 13646
rect 14702 13634 14754 13646
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 13794 13582 13806 13634
rect 13858 13582 13870 13634
rect 8318 13570 8370 13582
rect 14702 13570 14754 13582
rect 15262 13634 15314 13646
rect 15262 13570 15314 13582
rect 15486 13634 15538 13646
rect 31838 13634 31890 13646
rect 16706 13582 16718 13634
rect 16770 13582 16782 13634
rect 15486 13570 15538 13582
rect 31838 13570 31890 13582
rect 33182 13634 33234 13646
rect 36878 13634 36930 13646
rect 33506 13582 33518 13634
rect 33570 13582 33582 13634
rect 33182 13570 33234 13582
rect 36878 13570 36930 13582
rect 1344 13354 40544 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40544 13354
rect 1344 13268 40544 13302
rect 5742 13186 5794 13198
rect 5742 13122 5794 13134
rect 7422 13186 7474 13198
rect 7422 13122 7474 13134
rect 26686 13186 26738 13198
rect 26686 13122 26738 13134
rect 27246 13186 27298 13198
rect 32846 13186 32898 13198
rect 32274 13134 32286 13186
rect 32338 13134 32350 13186
rect 27246 13122 27298 13134
rect 32846 13122 32898 13134
rect 33070 13186 33122 13198
rect 33070 13122 33122 13134
rect 7646 13074 7698 13086
rect 7646 13010 7698 13022
rect 9662 13074 9714 13086
rect 33506 13022 33518 13074
rect 33570 13022 33582 13074
rect 9662 13010 9714 13022
rect 5518 12962 5570 12974
rect 5518 12898 5570 12910
rect 8654 12962 8706 12974
rect 9550 12962 9602 12974
rect 9202 12910 9214 12962
rect 9266 12910 9278 12962
rect 8654 12898 8706 12910
rect 9550 12898 9602 12910
rect 9998 12962 10050 12974
rect 19518 12962 19570 12974
rect 10658 12910 10670 12962
rect 10722 12910 10734 12962
rect 18722 12910 18734 12962
rect 18786 12910 18798 12962
rect 19058 12910 19070 12962
rect 19122 12910 19134 12962
rect 9998 12898 10050 12910
rect 19518 12898 19570 12910
rect 21198 12962 21250 12974
rect 21198 12898 21250 12910
rect 21534 12962 21586 12974
rect 21534 12898 21586 12910
rect 21870 12962 21922 12974
rect 21870 12898 21922 12910
rect 26350 12962 26402 12974
rect 26350 12898 26402 12910
rect 30718 12962 30770 12974
rect 30718 12898 30770 12910
rect 30830 12962 30882 12974
rect 30830 12898 30882 12910
rect 31054 12962 31106 12974
rect 31054 12898 31106 12910
rect 31278 12962 31330 12974
rect 31838 12962 31890 12974
rect 31490 12910 31502 12962
rect 31554 12910 31566 12962
rect 32610 12910 32622 12962
rect 32674 12910 32686 12962
rect 36418 12910 36430 12962
rect 36482 12910 36494 12962
rect 38882 12910 38894 12962
rect 38946 12910 38958 12962
rect 31278 12898 31330 12910
rect 31838 12898 31890 12910
rect 9886 12850 9938 12862
rect 11790 12850 11842 12862
rect 27134 12850 27186 12862
rect 31726 12850 31778 12862
rect 10434 12798 10446 12850
rect 10498 12798 10510 12850
rect 13906 12798 13918 12850
rect 13970 12798 13982 12850
rect 25554 12798 25566 12850
rect 25618 12798 25630 12850
rect 26002 12798 26014 12850
rect 26066 12798 26078 12850
rect 30258 12798 30270 12850
rect 30322 12798 30334 12850
rect 35634 12798 35646 12850
rect 35698 12798 35710 12850
rect 40002 12798 40014 12850
rect 40066 12798 40078 12850
rect 9886 12786 9938 12798
rect 11790 12786 11842 12798
rect 27134 12786 27186 12798
rect 31726 12786 31778 12798
rect 5854 12738 5906 12750
rect 5854 12674 5906 12686
rect 6078 12738 6130 12750
rect 6078 12674 6130 12686
rect 7870 12738 7922 12750
rect 7870 12674 7922 12686
rect 7982 12738 8034 12750
rect 7982 12674 8034 12686
rect 8094 12738 8146 12750
rect 8094 12674 8146 12686
rect 8766 12738 8818 12750
rect 8766 12674 8818 12686
rect 8878 12738 8930 12750
rect 8878 12674 8930 12686
rect 8990 12738 9042 12750
rect 8990 12674 9042 12686
rect 11902 12738 11954 12750
rect 11902 12674 11954 12686
rect 19294 12738 19346 12750
rect 19294 12674 19346 12686
rect 19406 12738 19458 12750
rect 19406 12674 19458 12686
rect 19630 12738 19682 12750
rect 19630 12674 19682 12686
rect 21422 12738 21474 12750
rect 21422 12674 21474 12686
rect 29934 12738 29986 12750
rect 29934 12674 29986 12686
rect 32734 12738 32786 12750
rect 32734 12674 32786 12686
rect 37102 12738 37154 12750
rect 37102 12674 37154 12686
rect 1344 12570 40544 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40544 12570
rect 1344 12484 40544 12518
rect 6302 12402 6354 12414
rect 9550 12402 9602 12414
rect 6626 12350 6638 12402
rect 6690 12350 6702 12402
rect 8418 12350 8430 12402
rect 8482 12350 8494 12402
rect 6302 12338 6354 12350
rect 9550 12338 9602 12350
rect 9774 12402 9826 12414
rect 9774 12338 9826 12350
rect 9998 12402 10050 12414
rect 9998 12338 10050 12350
rect 11230 12402 11282 12414
rect 13582 12402 13634 12414
rect 11554 12350 11566 12402
rect 11618 12350 11630 12402
rect 11230 12338 11282 12350
rect 13582 12338 13634 12350
rect 13694 12402 13746 12414
rect 13694 12338 13746 12350
rect 13806 12402 13858 12414
rect 18958 12402 19010 12414
rect 14914 12350 14926 12402
rect 14978 12350 14990 12402
rect 13806 12338 13858 12350
rect 18958 12338 19010 12350
rect 20526 12402 20578 12414
rect 20526 12338 20578 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 27918 12402 27970 12414
rect 27918 12338 27970 12350
rect 31838 12402 31890 12414
rect 31838 12338 31890 12350
rect 32286 12402 32338 12414
rect 32286 12338 32338 12350
rect 33182 12402 33234 12414
rect 33182 12338 33234 12350
rect 15934 12290 15986 12302
rect 15934 12226 15986 12238
rect 16382 12290 16434 12302
rect 20638 12290 20690 12302
rect 31166 12290 31218 12302
rect 17602 12238 17614 12290
rect 17666 12238 17678 12290
rect 30930 12238 30942 12290
rect 30994 12238 31006 12290
rect 16382 12226 16434 12238
rect 20638 12226 20690 12238
rect 31166 12226 31218 12238
rect 34078 12290 34130 12302
rect 34078 12226 34130 12238
rect 40126 12290 40178 12302
rect 40126 12226 40178 12238
rect 4846 12178 4898 12190
rect 4846 12114 4898 12126
rect 5294 12178 5346 12190
rect 5294 12114 5346 12126
rect 5742 12178 5794 12190
rect 5742 12114 5794 12126
rect 7870 12178 7922 12190
rect 7870 12114 7922 12126
rect 14254 12178 14306 12190
rect 14254 12114 14306 12126
rect 14590 12178 14642 12190
rect 17390 12178 17442 12190
rect 15698 12126 15710 12178
rect 15762 12126 15774 12178
rect 14590 12114 14642 12126
rect 17390 12114 17442 12126
rect 17838 12178 17890 12190
rect 20414 12178 20466 12190
rect 17938 12126 17950 12178
rect 18002 12126 18014 12178
rect 20066 12126 20078 12178
rect 20130 12126 20142 12178
rect 17838 12114 17890 12126
rect 20414 12114 20466 12126
rect 28030 12178 28082 12190
rect 28030 12114 28082 12126
rect 28590 12178 28642 12190
rect 28590 12114 28642 12126
rect 30830 12178 30882 12190
rect 30830 12114 30882 12126
rect 31614 12178 31666 12190
rect 31614 12114 31666 12126
rect 33630 12178 33682 12190
rect 33630 12114 33682 12126
rect 33742 12178 33794 12190
rect 33742 12114 33794 12126
rect 33966 12178 34018 12190
rect 33966 12114 34018 12126
rect 4510 12066 4562 12078
rect 4510 12002 4562 12014
rect 8094 12066 8146 12078
rect 8094 12002 8146 12014
rect 9662 12066 9714 12078
rect 9662 12002 9714 12014
rect 14030 12066 14082 12078
rect 14030 12002 14082 12014
rect 16494 12066 16546 12078
rect 16494 12002 16546 12014
rect 16606 12066 16658 12078
rect 16606 12002 16658 12014
rect 17502 12066 17554 12078
rect 17502 12002 17554 12014
rect 21086 12066 21138 12078
rect 21086 12002 21138 12014
rect 5070 11954 5122 11966
rect 5070 11890 5122 11902
rect 25230 11954 25282 11966
rect 25230 11890 25282 11902
rect 25566 11954 25618 11966
rect 25566 11890 25618 11902
rect 27918 11954 27970 11966
rect 27918 11890 27970 11902
rect 28702 11954 28754 11966
rect 28702 11890 28754 11902
rect 1344 11786 40544 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40544 11786
rect 1344 11700 40544 11734
rect 19854 11618 19906 11630
rect 17602 11566 17614 11618
rect 17666 11566 17678 11618
rect 19854 11554 19906 11566
rect 9214 11506 9266 11518
rect 4834 11454 4846 11506
rect 4898 11454 4910 11506
rect 9214 11442 9266 11454
rect 10558 11506 10610 11518
rect 10558 11442 10610 11454
rect 13470 11506 13522 11518
rect 13470 11442 13522 11454
rect 15150 11506 15202 11518
rect 15150 11442 15202 11454
rect 18622 11506 18674 11518
rect 18622 11442 18674 11454
rect 23214 11506 23266 11518
rect 23214 11442 23266 11454
rect 25118 11506 25170 11518
rect 25118 11442 25170 11454
rect 33854 11506 33906 11518
rect 33854 11442 33906 11454
rect 5630 11394 5682 11406
rect 2034 11342 2046 11394
rect 2098 11342 2110 11394
rect 5630 11330 5682 11342
rect 6750 11394 6802 11406
rect 7982 11394 8034 11406
rect 7186 11342 7198 11394
rect 7250 11342 7262 11394
rect 6750 11330 6802 11342
rect 7982 11330 8034 11342
rect 8430 11394 8482 11406
rect 9438 11394 9490 11406
rect 8754 11342 8766 11394
rect 8818 11342 8830 11394
rect 8430 11330 8482 11342
rect 9438 11330 9490 11342
rect 9774 11394 9826 11406
rect 9774 11330 9826 11342
rect 13582 11394 13634 11406
rect 16830 11394 16882 11406
rect 14130 11342 14142 11394
rect 14194 11342 14206 11394
rect 13582 11330 13634 11342
rect 16830 11330 16882 11342
rect 17166 11394 17218 11406
rect 17838 11394 17890 11406
rect 17602 11342 17614 11394
rect 17666 11342 17678 11394
rect 17166 11330 17218 11342
rect 17838 11330 17890 11342
rect 18174 11394 18226 11406
rect 25006 11394 25058 11406
rect 20178 11342 20190 11394
rect 20242 11342 20254 11394
rect 20402 11342 20414 11394
rect 20466 11342 20478 11394
rect 21522 11342 21534 11394
rect 21586 11342 21598 11394
rect 24434 11342 24446 11394
rect 24498 11342 24510 11394
rect 18174 11330 18226 11342
rect 25006 11330 25058 11342
rect 29150 11394 29202 11406
rect 29150 11330 29202 11342
rect 32958 11394 33010 11406
rect 32958 11330 33010 11342
rect 7646 11282 7698 11294
rect 10110 11282 10162 11294
rect 2706 11230 2718 11282
rect 2770 11230 2782 11282
rect 5954 11230 5966 11282
rect 6018 11230 6030 11282
rect 8194 11230 8206 11282
rect 8258 11230 8270 11282
rect 7646 11218 7698 11230
rect 10110 11218 10162 11230
rect 16942 11282 16994 11294
rect 28142 11282 28194 11294
rect 18946 11230 18958 11282
rect 19010 11230 19022 11282
rect 21298 11230 21310 11282
rect 21362 11230 21374 11282
rect 16942 11218 16994 11230
rect 28142 11218 28194 11230
rect 28254 11282 28306 11294
rect 28254 11218 28306 11230
rect 29486 11282 29538 11294
rect 33282 11230 33294 11282
rect 33346 11230 33358 11282
rect 29486 11218 29538 11230
rect 8766 11170 8818 11182
rect 8766 11106 8818 11118
rect 9662 11170 9714 11182
rect 9662 11106 9714 11118
rect 17390 11170 17442 11182
rect 17390 11106 17442 11118
rect 19294 11170 19346 11182
rect 19294 11106 19346 11118
rect 19966 11170 20018 11182
rect 19966 11106 20018 11118
rect 27918 11170 27970 11182
rect 27918 11106 27970 11118
rect 29262 11170 29314 11182
rect 29262 11106 29314 11118
rect 31950 11170 32002 11182
rect 31950 11106 32002 11118
rect 1344 11002 40544 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40544 11002
rect 1344 10916 40544 10950
rect 6302 10834 6354 10846
rect 5842 10782 5854 10834
rect 5906 10782 5918 10834
rect 6302 10770 6354 10782
rect 7534 10834 7586 10846
rect 7534 10770 7586 10782
rect 8318 10834 8370 10846
rect 11902 10834 11954 10846
rect 8754 10782 8766 10834
rect 8818 10782 8830 10834
rect 8318 10770 8370 10782
rect 7646 10722 7698 10734
rect 7646 10658 7698 10670
rect 8206 10722 8258 10734
rect 8530 10670 8542 10722
rect 8594 10719 8606 10722
rect 8769 10719 8815 10782
rect 11902 10770 11954 10782
rect 12350 10834 12402 10846
rect 12350 10770 12402 10782
rect 25454 10834 25506 10846
rect 29934 10834 29986 10846
rect 27570 10782 27582 10834
rect 27634 10782 27646 10834
rect 25454 10770 25506 10782
rect 29934 10770 29986 10782
rect 8594 10673 8815 10719
rect 10558 10722 10610 10734
rect 24334 10722 24386 10734
rect 8594 10670 8606 10673
rect 19618 10670 19630 10722
rect 19682 10670 19694 10722
rect 28914 10670 28926 10722
rect 28978 10670 28990 10722
rect 8206 10658 8258 10670
rect 10558 10658 10610 10670
rect 24334 10658 24386 10670
rect 5518 10610 5570 10622
rect 8430 10610 8482 10622
rect 2370 10558 2382 10610
rect 2434 10558 2446 10610
rect 3042 10558 3054 10610
rect 3106 10558 3118 10610
rect 7298 10558 7310 10610
rect 7362 10558 7374 10610
rect 5518 10546 5570 10558
rect 8430 10546 8482 10558
rect 9662 10610 9714 10622
rect 9662 10546 9714 10558
rect 9774 10610 9826 10622
rect 9774 10546 9826 10558
rect 9998 10610 10050 10622
rect 9998 10546 10050 10558
rect 10110 10610 10162 10622
rect 10110 10546 10162 10558
rect 12126 10610 12178 10622
rect 24222 10610 24274 10622
rect 12562 10558 12574 10610
rect 12626 10558 12638 10610
rect 12898 10558 12910 10610
rect 12962 10558 12974 10610
rect 22978 10558 22990 10610
rect 23042 10558 23054 10610
rect 23650 10558 23662 10610
rect 23714 10558 23726 10610
rect 12126 10546 12178 10558
rect 24222 10546 24274 10558
rect 25342 10610 25394 10622
rect 25342 10546 25394 10558
rect 25566 10610 25618 10622
rect 25566 10546 25618 10558
rect 26014 10610 26066 10622
rect 29710 10610 29762 10622
rect 27906 10558 27918 10610
rect 27970 10558 27982 10610
rect 28578 10558 28590 10610
rect 28642 10558 28654 10610
rect 26014 10546 26066 10558
rect 29710 10546 29762 10558
rect 30046 10610 30098 10622
rect 30046 10546 30098 10558
rect 30270 10610 30322 10622
rect 36878 10610 36930 10622
rect 36418 10558 36430 10610
rect 36482 10558 36494 10610
rect 30270 10546 30322 10558
rect 36878 10546 36930 10558
rect 8878 10498 8930 10510
rect 5170 10446 5182 10498
rect 5234 10446 5246 10498
rect 8878 10434 8930 10446
rect 12238 10498 12290 10510
rect 12238 10434 12290 10446
rect 13358 10498 13410 10510
rect 33506 10446 33518 10498
rect 33570 10446 33582 10498
rect 35634 10446 35646 10498
rect 35698 10446 35710 10498
rect 13358 10434 13410 10446
rect 1344 10218 40544 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40544 10218
rect 1344 10132 40544 10166
rect 8654 10050 8706 10062
rect 8654 9986 8706 9998
rect 21422 10050 21474 10062
rect 21422 9986 21474 9998
rect 29150 10050 29202 10062
rect 29150 9986 29202 9998
rect 29486 10050 29538 10062
rect 29486 9986 29538 9998
rect 12126 9938 12178 9950
rect 12126 9874 12178 9886
rect 14030 9938 14082 9950
rect 20750 9938 20802 9950
rect 23662 9938 23714 9950
rect 25342 9938 25394 9950
rect 16034 9886 16046 9938
rect 16098 9886 16110 9938
rect 18162 9886 18174 9938
rect 18226 9886 18238 9938
rect 18610 9886 18622 9938
rect 18674 9886 18686 9938
rect 20514 9886 20526 9938
rect 20578 9886 20590 9938
rect 22306 9886 22318 9938
rect 22370 9886 22382 9938
rect 24770 9886 24782 9938
rect 24834 9886 24846 9938
rect 14030 9874 14082 9886
rect 20750 9874 20802 9886
rect 23662 9874 23714 9886
rect 25342 9874 25394 9886
rect 30942 9938 30994 9950
rect 30942 9874 30994 9886
rect 31390 9938 31442 9950
rect 34078 9938 34130 9950
rect 32834 9886 32846 9938
rect 32898 9886 32910 9938
rect 34850 9886 34862 9938
rect 34914 9886 34926 9938
rect 31390 9874 31442 9886
rect 34078 9874 34130 9886
rect 22206 9826 22258 9838
rect 8978 9774 8990 9826
rect 9042 9774 9054 9826
rect 15362 9774 15374 9826
rect 15426 9774 15438 9826
rect 21746 9774 21758 9826
rect 21810 9774 21822 9826
rect 22206 9762 22258 9774
rect 23214 9826 23266 9838
rect 23214 9762 23266 9774
rect 23438 9826 23490 9838
rect 23438 9762 23490 9774
rect 23886 9826 23938 9838
rect 34190 9826 34242 9838
rect 24210 9774 24222 9826
rect 24274 9774 24286 9826
rect 26898 9774 26910 9826
rect 26962 9774 26974 9826
rect 27794 9774 27806 9826
rect 27858 9774 27870 9826
rect 32610 9774 32622 9826
rect 32674 9774 32686 9826
rect 33842 9774 33854 9826
rect 33906 9774 33918 9826
rect 23886 9762 23938 9774
rect 34190 9762 34242 9774
rect 19070 9714 19122 9726
rect 21310 9714 21362 9726
rect 19730 9662 19742 9714
rect 19794 9662 19806 9714
rect 19070 9650 19122 9662
rect 21310 9650 21362 9662
rect 24782 9714 24834 9726
rect 29374 9714 29426 9726
rect 26338 9662 26350 9714
rect 26402 9662 26414 9714
rect 24782 9650 24834 9662
rect 29374 9650 29426 9662
rect 33294 9714 33346 9726
rect 33294 9650 33346 9662
rect 34526 9714 34578 9726
rect 34526 9650 34578 9662
rect 34750 9714 34802 9726
rect 34750 9650 34802 9662
rect 8766 9602 8818 9614
rect 8766 9538 8818 9550
rect 9438 9602 9490 9614
rect 9438 9538 9490 9550
rect 12014 9602 12066 9614
rect 12014 9538 12066 9550
rect 20078 9602 20130 9614
rect 20078 9538 20130 9550
rect 21982 9602 22034 9614
rect 21982 9538 22034 9550
rect 22318 9602 22370 9614
rect 22318 9538 22370 9550
rect 22878 9602 22930 9614
rect 22878 9538 22930 9550
rect 24446 9602 24498 9614
rect 24446 9538 24498 9550
rect 24670 9602 24722 9614
rect 24670 9538 24722 9550
rect 25230 9602 25282 9614
rect 30382 9602 30434 9614
rect 27906 9550 27918 9602
rect 27970 9550 27982 9602
rect 25230 9538 25282 9550
rect 30382 9538 30434 9550
rect 31950 9602 32002 9614
rect 31950 9538 32002 9550
rect 1344 9434 40544 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40544 9434
rect 1344 9348 40544 9382
rect 24558 9266 24610 9278
rect 24558 9202 24610 9214
rect 25678 9266 25730 9278
rect 25678 9202 25730 9214
rect 26014 9266 26066 9278
rect 26014 9202 26066 9214
rect 26238 9266 26290 9278
rect 26238 9202 26290 9214
rect 28142 9266 28194 9278
rect 28142 9202 28194 9214
rect 28254 9266 28306 9278
rect 28254 9202 28306 9214
rect 29150 9266 29202 9278
rect 29150 9202 29202 9214
rect 18734 9154 18786 9166
rect 11666 9102 11678 9154
rect 11730 9102 11742 9154
rect 18734 9090 18786 9102
rect 18958 9154 19010 9166
rect 23774 9154 23826 9166
rect 20626 9102 20638 9154
rect 20690 9102 20702 9154
rect 18958 9090 19010 9102
rect 23774 9090 23826 9102
rect 23886 9154 23938 9166
rect 23886 9090 23938 9102
rect 25230 9154 25282 9166
rect 25230 9090 25282 9102
rect 25454 9154 25506 9166
rect 25454 9090 25506 9102
rect 27806 9154 27858 9166
rect 27806 9090 27858 9102
rect 28590 9154 28642 9166
rect 31714 9102 31726 9154
rect 31778 9102 31790 9154
rect 35186 9102 35198 9154
rect 35250 9102 35262 9154
rect 28590 9090 28642 9102
rect 19294 9042 19346 9054
rect 10882 8990 10894 9042
rect 10946 8990 10958 9042
rect 14914 8990 14926 9042
rect 14978 8990 14990 9042
rect 19294 8978 19346 8990
rect 19406 9042 19458 9054
rect 24670 9042 24722 9054
rect 19842 8990 19854 9042
rect 19906 8990 19918 9042
rect 24322 8990 24334 9042
rect 24386 8990 24398 9042
rect 19406 8978 19458 8990
rect 24670 8978 24722 8990
rect 25902 9042 25954 9054
rect 25902 8978 25954 8990
rect 26350 9042 26402 9054
rect 27694 9042 27746 9054
rect 27122 8990 27134 9042
rect 27186 8990 27198 9042
rect 26350 8978 26402 8990
rect 27694 8978 27746 8990
rect 28366 9042 28418 9054
rect 36430 9042 36482 9054
rect 32498 8990 32510 9042
rect 32562 8990 32574 9042
rect 35858 8990 35870 9042
rect 35922 8990 35934 9042
rect 28366 8978 28418 8990
rect 36430 8978 36482 8990
rect 14254 8930 14306 8942
rect 19070 8930 19122 8942
rect 13794 8878 13806 8930
rect 13858 8878 13870 8930
rect 14690 8878 14702 8930
rect 14754 8878 14766 8930
rect 22754 8878 22766 8930
rect 22818 8878 22830 8930
rect 29586 8878 29598 8930
rect 29650 8878 29662 8930
rect 33058 8878 33070 8930
rect 33122 8878 33134 8930
rect 14254 8866 14306 8878
rect 19070 8866 19122 8878
rect 1344 8650 40544 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40544 8650
rect 1344 8564 40544 8598
rect 14590 8482 14642 8494
rect 14590 8418 14642 8430
rect 28366 8482 28418 8494
rect 28366 8418 28418 8430
rect 32286 8482 32338 8494
rect 32286 8418 32338 8430
rect 11454 8370 11506 8382
rect 20078 8370 20130 8382
rect 8866 8318 8878 8370
rect 8930 8318 8942 8370
rect 10994 8318 11006 8370
rect 11058 8318 11070 8370
rect 14242 8318 14254 8370
rect 14306 8318 14318 8370
rect 17042 8318 17054 8370
rect 17106 8318 17118 8370
rect 19170 8318 19182 8370
rect 19234 8318 19246 8370
rect 11454 8306 11506 8318
rect 20078 8306 20130 8318
rect 20302 8370 20354 8382
rect 20302 8306 20354 8318
rect 26126 8370 26178 8382
rect 26126 8306 26178 8318
rect 27806 8370 27858 8382
rect 27806 8306 27858 8318
rect 32398 8370 32450 8382
rect 32398 8306 32450 8318
rect 19966 8258 20018 8270
rect 21646 8258 21698 8270
rect 27918 8258 27970 8270
rect 8082 8206 8094 8258
rect 8146 8206 8158 8258
rect 16370 8206 16382 8258
rect 16434 8206 16446 8258
rect 20514 8206 20526 8258
rect 20578 8206 20590 8258
rect 22082 8206 22094 8258
rect 22146 8206 22158 8258
rect 27570 8206 27582 8258
rect 27634 8206 27646 8258
rect 19966 8194 20018 8206
rect 21646 8194 21698 8206
rect 27918 8194 27970 8206
rect 28254 8258 28306 8270
rect 38882 8206 38894 8258
rect 38946 8206 38958 8258
rect 28254 8194 28306 8206
rect 14030 8146 14082 8158
rect 14030 8082 14082 8094
rect 21422 8146 21474 8158
rect 21422 8082 21474 8094
rect 21534 8146 21586 8158
rect 22754 8094 22766 8146
rect 22818 8094 22830 8146
rect 40002 8094 40014 8146
rect 40066 8094 40078 8146
rect 21534 8082 21586 8094
rect 14366 8034 14418 8046
rect 14366 7970 14418 7982
rect 15038 8034 15090 8046
rect 15038 7970 15090 7982
rect 19742 8034 19794 8046
rect 19742 7970 19794 7982
rect 22430 8034 22482 8046
rect 22430 7970 22482 7982
rect 28366 8034 28418 8046
rect 28366 7970 28418 7982
rect 32846 8034 32898 8046
rect 32846 7970 32898 7982
rect 1344 7866 40544 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40544 7866
rect 1344 7780 40544 7814
rect 21086 7698 21138 7710
rect 21086 7634 21138 7646
rect 40126 7698 40178 7710
rect 40126 7634 40178 7646
rect 39678 7586 39730 7598
rect 13906 7534 13918 7586
rect 13970 7534 13982 7586
rect 39678 7522 39730 7534
rect 16494 7474 16546 7486
rect 13122 7422 13134 7474
rect 13186 7422 13198 7474
rect 16494 7410 16546 7422
rect 16034 7310 16046 7362
rect 16098 7310 16110 7362
rect 1344 7082 40544 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40544 7082
rect 1344 6996 40544 7030
rect 25566 6914 25618 6926
rect 25566 6850 25618 6862
rect 25230 6802 25282 6814
rect 25230 6738 25282 6750
rect 21310 6690 21362 6702
rect 21310 6626 21362 6638
rect 21534 6690 21586 6702
rect 26462 6690 26514 6702
rect 21858 6638 21870 6690
rect 21922 6638 21934 6690
rect 22306 6638 22318 6690
rect 22370 6638 22382 6690
rect 21534 6626 21586 6638
rect 26462 6626 26514 6638
rect 27470 6690 27522 6702
rect 27470 6626 27522 6638
rect 22990 6578 23042 6590
rect 22530 6526 22542 6578
rect 22594 6526 22606 6578
rect 22990 6514 23042 6526
rect 24222 6578 24274 6590
rect 24222 6514 24274 6526
rect 24334 6578 24386 6590
rect 24334 6514 24386 6526
rect 24894 6578 24946 6590
rect 24894 6514 24946 6526
rect 25454 6578 25506 6590
rect 25454 6514 25506 6526
rect 26014 6578 26066 6590
rect 26014 6514 26066 6526
rect 1710 6466 1762 6478
rect 1710 6402 1762 6414
rect 21422 6466 21474 6478
rect 21422 6402 21474 6414
rect 24558 6466 24610 6478
rect 24558 6402 24610 6414
rect 25902 6466 25954 6478
rect 40126 6466 40178 6478
rect 27122 6414 27134 6466
rect 27186 6414 27198 6466
rect 25902 6402 25954 6414
rect 40126 6402 40178 6414
rect 1344 6298 40544 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40544 6298
rect 1344 6212 40544 6246
rect 23214 6130 23266 6142
rect 23214 6066 23266 6078
rect 1710 6018 1762 6030
rect 23438 6018 23490 6030
rect 19506 5966 19518 6018
rect 19570 5966 19582 6018
rect 1710 5954 1762 5966
rect 23438 5954 23490 5966
rect 24670 6018 24722 6030
rect 39790 6018 39842 6030
rect 26226 5966 26238 6018
rect 26290 5966 26302 6018
rect 24670 5954 24722 5966
rect 39790 5954 39842 5966
rect 21982 5906 22034 5918
rect 18834 5854 18846 5906
rect 18898 5854 18910 5906
rect 21982 5842 22034 5854
rect 22206 5906 22258 5918
rect 22206 5842 22258 5854
rect 23102 5906 23154 5918
rect 28814 5906 28866 5918
rect 24098 5854 24110 5906
rect 24162 5854 24174 5906
rect 25554 5854 25566 5906
rect 25618 5854 25630 5906
rect 23102 5842 23154 5854
rect 28814 5842 28866 5854
rect 39566 5906 39618 5918
rect 39566 5842 39618 5854
rect 40126 5906 40178 5918
rect 40126 5842 40178 5854
rect 21634 5742 21646 5794
rect 21698 5742 21710 5794
rect 24210 5742 24222 5794
rect 24274 5742 24286 5794
rect 28354 5742 28366 5794
rect 28418 5742 28430 5794
rect 22530 5630 22542 5682
rect 22594 5630 22606 5682
rect 1344 5514 40544 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40544 5514
rect 1344 5428 40544 5462
rect 21310 5346 21362 5358
rect 21310 5282 21362 5294
rect 26126 5346 26178 5358
rect 26126 5282 26178 5294
rect 25778 5182 25790 5234
rect 25842 5182 25854 5234
rect 26238 5122 26290 5134
rect 21634 5070 21646 5122
rect 21698 5070 21710 5122
rect 22866 5070 22878 5122
rect 22930 5070 22942 5122
rect 26450 5070 26462 5122
rect 26514 5070 26526 5122
rect 38434 5070 38446 5122
rect 38498 5070 38510 5122
rect 26238 5058 26290 5070
rect 38670 5010 38722 5022
rect 23650 4958 23662 5010
rect 23714 4958 23726 5010
rect 38670 4946 38722 4958
rect 1710 4898 1762 4910
rect 1710 4834 1762 4846
rect 21422 4898 21474 4910
rect 21422 4834 21474 4846
rect 40126 4898 40178 4910
rect 40126 4834 40178 4846
rect 1344 4730 40544 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40544 4730
rect 1344 4644 40544 4678
rect 24110 4562 24162 4574
rect 24110 4498 24162 4510
rect 1710 4450 1762 4462
rect 24334 4450 24386 4462
rect 20178 4398 20190 4450
rect 20242 4398 20254 4450
rect 1710 4386 1762 4398
rect 24334 4386 24386 4398
rect 39678 4450 39730 4462
rect 39678 4386 39730 4398
rect 40126 4450 40178 4462
rect 40126 4386 40178 4398
rect 19506 4286 19518 4338
rect 19570 4286 19582 4338
rect 22306 4174 22318 4226
rect 22370 4174 22382 4226
rect 23986 4174 23998 4226
rect 24050 4174 24062 4226
rect 1344 3946 40544 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40544 3946
rect 1344 3860 40544 3894
rect 21186 3614 21198 3666
rect 21250 3614 21262 3666
rect 20750 3554 20802 3566
rect 20750 3490 20802 3502
rect 19630 3442 19682 3454
rect 19630 3378 19682 3390
rect 19854 3442 19906 3454
rect 19854 3378 19906 3390
rect 20190 3442 20242 3454
rect 20190 3378 20242 3390
rect 1710 3330 1762 3342
rect 1710 3266 1762 3278
rect 10334 3330 10386 3342
rect 10334 3266 10386 3278
rect 11006 3330 11058 3342
rect 11006 3266 11058 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 39230 3330 39282 3342
rect 39230 3266 39282 3278
rect 40126 3330 40178 3342
rect 40126 3266 40178 3278
rect 1344 3162 40544 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40544 3162
rect 1344 3076 40544 3110
<< via1 >>
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 8318 42142 8370 42194
rect 35982 42142 36034 42194
rect 38782 42142 38834 42194
rect 40126 42142 40178 42194
rect 39230 42030 39282 42082
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 39678 41022 39730 41074
rect 1710 40910 1762 40962
rect 29374 40910 29426 40962
rect 30382 40910 30434 40962
rect 30830 40910 30882 40962
rect 40126 40910 40178 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 40126 40462 40178 40514
rect 25902 40350 25954 40402
rect 29150 40350 29202 40402
rect 29598 40350 29650 40402
rect 26574 40238 26626 40290
rect 28702 40238 28754 40290
rect 30382 40238 30434 40290
rect 32510 40238 32562 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 27246 39790 27298 39842
rect 26350 39678 26402 39730
rect 31166 39678 31218 39730
rect 31838 39678 31890 39730
rect 31950 39678 32002 39730
rect 23550 39566 23602 39618
rect 29374 39566 29426 39618
rect 30830 39566 30882 39618
rect 32734 39566 32786 39618
rect 24222 39454 24274 39506
rect 27358 39454 27410 39506
rect 27582 39454 27634 39506
rect 31502 39454 31554 39506
rect 32062 39454 32114 39506
rect 26798 39342 26850 39394
rect 29150 39342 29202 39394
rect 29934 39342 29986 39394
rect 30046 39342 30098 39394
rect 30158 39342 30210 39394
rect 30382 39342 30434 39394
rect 31054 39342 31106 39394
rect 31278 39342 31330 39394
rect 32510 39342 32562 39394
rect 40126 39342 40178 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 25342 39006 25394 39058
rect 29822 39006 29874 39058
rect 31390 38894 31442 38946
rect 32062 38894 32114 38946
rect 33070 38894 33122 38946
rect 33294 38894 33346 38946
rect 40126 38894 40178 38946
rect 11342 38782 11394 38834
rect 25566 38782 25618 38834
rect 28254 38782 28306 38834
rect 30046 38782 30098 38834
rect 30942 38782 30994 38834
rect 32398 38782 32450 38834
rect 12014 38670 12066 38722
rect 14142 38670 14194 38722
rect 25230 38670 25282 38722
rect 27918 38670 27970 38722
rect 28814 38670 28866 38722
rect 33182 38670 33234 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 12350 38222 12402 38274
rect 31502 38222 31554 38274
rect 31726 38222 31778 38274
rect 14254 38110 14306 38162
rect 16270 38110 16322 38162
rect 21534 38110 21586 38162
rect 25118 38110 25170 38162
rect 28030 38110 28082 38162
rect 29374 38110 29426 38162
rect 30158 38110 30210 38162
rect 14142 37998 14194 38050
rect 19182 37998 19234 38050
rect 25342 37998 25394 38050
rect 26126 37998 26178 38050
rect 26574 37998 26626 38050
rect 27918 37998 27970 38050
rect 28366 37998 28418 38050
rect 29710 37998 29762 38050
rect 31166 37998 31218 38050
rect 12686 37886 12738 37938
rect 13470 37886 13522 37938
rect 15486 37886 15538 37938
rect 18398 37886 18450 37938
rect 21422 37886 21474 37938
rect 21646 37886 21698 37938
rect 24670 37886 24722 37938
rect 25118 37886 25170 37938
rect 26686 37886 26738 37938
rect 27358 37886 27410 37938
rect 28590 37886 28642 37938
rect 30494 37886 30546 37938
rect 30942 37886 30994 37938
rect 12462 37774 12514 37826
rect 14814 37774 14866 37826
rect 15150 37774 15202 37826
rect 15598 37774 15650 37826
rect 15822 37774 15874 37826
rect 19630 37774 19682 37826
rect 24894 37774 24946 37826
rect 28142 37774 28194 37826
rect 30606 37774 30658 37826
rect 31838 37774 31890 37826
rect 32174 37774 32226 37826
rect 32510 37774 32562 37826
rect 40126 37774 40178 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 9662 37438 9714 37490
rect 17614 37438 17666 37490
rect 23214 37438 23266 37490
rect 27470 37438 27522 37490
rect 28030 37438 28082 37490
rect 30606 37438 30658 37490
rect 31278 37438 31330 37490
rect 1710 37326 1762 37378
rect 16718 37326 16770 37378
rect 17390 37326 17442 37378
rect 21758 37326 21810 37378
rect 26574 37326 26626 37378
rect 30382 37326 30434 37378
rect 32062 37326 32114 37378
rect 40126 37326 40178 37378
rect 13470 37214 13522 37266
rect 15486 37214 15538 37266
rect 16158 37214 16210 37266
rect 16382 37214 16434 37266
rect 17838 37214 17890 37266
rect 22542 37214 22594 37266
rect 22878 37214 22930 37266
rect 26462 37214 26514 37266
rect 27358 37214 27410 37266
rect 30270 37214 30322 37266
rect 30718 37214 30770 37266
rect 31166 37214 31218 37266
rect 31390 37214 31442 37266
rect 31726 37214 31778 37266
rect 13582 37102 13634 37154
rect 14030 37102 14082 37154
rect 14814 37102 14866 37154
rect 15710 37102 15762 37154
rect 16606 37102 16658 37154
rect 19630 37102 19682 37154
rect 23662 37102 23714 37154
rect 25566 37102 25618 37154
rect 9550 36990 9602 37042
rect 9886 36990 9938 37042
rect 17278 36990 17330 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 14926 36654 14978 36706
rect 27022 36654 27074 36706
rect 8206 36542 8258 36594
rect 10334 36542 10386 36594
rect 12126 36542 12178 36594
rect 13806 36542 13858 36594
rect 15150 36542 15202 36594
rect 16942 36542 16994 36594
rect 24894 36542 24946 36594
rect 25790 36542 25842 36594
rect 26462 36542 26514 36594
rect 7534 36430 7586 36482
rect 12014 36430 12066 36482
rect 13582 36430 13634 36482
rect 13694 36430 13746 36482
rect 14030 36430 14082 36482
rect 16046 36430 16098 36482
rect 16718 36430 16770 36482
rect 17838 36430 17890 36482
rect 19406 36430 19458 36482
rect 20190 36430 20242 36482
rect 20750 36430 20802 36482
rect 21534 36430 21586 36482
rect 21646 36430 21698 36482
rect 21758 36430 21810 36482
rect 21870 36430 21922 36482
rect 25454 36430 25506 36482
rect 26686 36430 26738 36482
rect 29374 36430 29426 36482
rect 1710 36318 1762 36370
rect 12686 36318 12738 36370
rect 15822 36318 15874 36370
rect 18958 36318 19010 36370
rect 29150 36318 29202 36370
rect 12238 36206 12290 36258
rect 12462 36206 12514 36258
rect 13918 36206 13970 36258
rect 14590 36206 14642 36258
rect 16382 36206 16434 36258
rect 17166 36206 17218 36258
rect 17278 36206 17330 36258
rect 17390 36206 17442 36258
rect 18174 36206 18226 36258
rect 21422 36206 21474 36258
rect 22542 36206 22594 36258
rect 31278 36206 31330 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 8430 35870 8482 35922
rect 15934 35870 15986 35922
rect 17726 35870 17778 35922
rect 20862 35870 20914 35922
rect 23326 35870 23378 35922
rect 9774 35758 9826 35810
rect 9998 35758 10050 35810
rect 11678 35758 11730 35810
rect 15710 35758 15762 35810
rect 16494 35758 16546 35810
rect 16606 35758 16658 35810
rect 17390 35758 17442 35810
rect 17502 35758 17554 35810
rect 30382 35758 30434 35810
rect 31502 35758 31554 35810
rect 32286 35758 32338 35810
rect 8206 35646 8258 35698
rect 11230 35646 11282 35698
rect 13694 35646 13746 35698
rect 15598 35646 15650 35698
rect 20526 35646 20578 35698
rect 23550 35646 23602 35698
rect 26798 35646 26850 35698
rect 31278 35646 31330 35698
rect 32510 35646 32562 35698
rect 33070 35646 33122 35698
rect 8878 35534 8930 35586
rect 13470 35534 13522 35586
rect 18062 35534 18114 35586
rect 22990 35534 23042 35586
rect 24782 35534 24834 35586
rect 32174 35534 32226 35586
rect 33182 35534 33234 35586
rect 14030 35422 14082 35474
rect 16494 35422 16546 35474
rect 30942 35422 30994 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 11678 35086 11730 35138
rect 11230 34974 11282 35026
rect 15262 34974 15314 35026
rect 16830 34974 16882 35026
rect 25902 34974 25954 35026
rect 27246 34974 27298 35026
rect 34526 34974 34578 35026
rect 10222 34862 10274 34914
rect 10782 34862 10834 34914
rect 12014 34862 12066 34914
rect 14702 34862 14754 34914
rect 19742 34862 19794 34914
rect 23102 34862 23154 34914
rect 26238 34862 26290 34914
rect 26686 34862 26738 34914
rect 30830 34862 30882 34914
rect 31614 34862 31666 34914
rect 10446 34750 10498 34802
rect 18846 34750 18898 34802
rect 18958 34750 19010 34802
rect 19406 34750 19458 34802
rect 23774 34750 23826 34802
rect 30494 34750 30546 34802
rect 32398 34750 32450 34802
rect 11790 34638 11842 34690
rect 14926 34638 14978 34690
rect 15150 34638 15202 34690
rect 15262 34638 15314 34690
rect 16382 34638 16434 34690
rect 19182 34638 19234 34690
rect 19518 34638 19570 34690
rect 29934 34638 29986 34690
rect 30158 34638 30210 34690
rect 30382 34638 30434 34690
rect 31054 34638 31106 34690
rect 31278 34638 31330 34690
rect 31390 34638 31442 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 7870 34302 7922 34354
rect 9774 34302 9826 34354
rect 13246 34302 13298 34354
rect 13582 34302 13634 34354
rect 15710 34302 15762 34354
rect 16270 34302 16322 34354
rect 23438 34302 23490 34354
rect 23886 34302 23938 34354
rect 30494 34302 30546 34354
rect 31278 34302 31330 34354
rect 8990 34190 9042 34242
rect 12014 34190 12066 34242
rect 16046 34190 16098 34242
rect 16494 34190 16546 34242
rect 19518 34190 19570 34242
rect 25790 34190 25842 34242
rect 29710 34190 29762 34242
rect 30270 34190 30322 34242
rect 31054 34190 31106 34242
rect 31390 34190 31442 34242
rect 33070 34190 33122 34242
rect 8766 34078 8818 34130
rect 9662 34078 9714 34130
rect 9886 34078 9938 34130
rect 10334 34078 10386 34130
rect 10558 34078 10610 34130
rect 11790 34078 11842 34130
rect 12126 34078 12178 34130
rect 15374 34078 15426 34130
rect 16606 34078 16658 34130
rect 19182 34078 19234 34130
rect 20190 34078 20242 34130
rect 20302 34078 20354 34130
rect 20526 34078 20578 34130
rect 23662 34078 23714 34130
rect 24110 34078 24162 34130
rect 24334 34078 24386 34130
rect 26126 34078 26178 34130
rect 29038 34078 29090 34130
rect 29374 34078 29426 34130
rect 30158 34078 30210 34130
rect 30942 34078 30994 34130
rect 32286 34078 32338 34130
rect 33518 34078 33570 34130
rect 33966 34078 34018 34130
rect 10894 33966 10946 34018
rect 14254 33966 14306 34018
rect 15150 33966 15202 34018
rect 16382 33966 16434 34018
rect 31838 33966 31890 34018
rect 7758 33854 7810 33906
rect 8094 33854 8146 33906
rect 20638 33854 20690 33906
rect 31614 33854 31666 33906
rect 31838 33854 31890 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 13806 33518 13858 33570
rect 18622 33518 18674 33570
rect 32174 33518 32226 33570
rect 5630 33406 5682 33458
rect 7758 33406 7810 33458
rect 9214 33406 9266 33458
rect 11006 33406 11058 33458
rect 13470 33406 13522 33458
rect 14926 33406 14978 33458
rect 15374 33406 15426 33458
rect 15822 33406 15874 33458
rect 20078 33406 20130 33458
rect 27918 33406 27970 33458
rect 28478 33406 28530 33458
rect 30270 33406 30322 33458
rect 8542 33294 8594 33346
rect 9550 33294 9602 33346
rect 11118 33294 11170 33346
rect 11342 33294 11394 33346
rect 14814 33294 14866 33346
rect 15038 33294 15090 33346
rect 16046 33294 16098 33346
rect 18398 33294 18450 33346
rect 19294 33294 19346 33346
rect 25118 33294 25170 33346
rect 30382 33294 30434 33346
rect 35198 33294 35250 33346
rect 8878 33182 8930 33234
rect 10670 33182 10722 33234
rect 11566 33182 11618 33234
rect 11678 33182 11730 33234
rect 13582 33182 13634 33234
rect 14478 33182 14530 33234
rect 19518 33182 19570 33234
rect 19630 33238 19682 33290
rect 19854 33182 19906 33234
rect 22094 33182 22146 33234
rect 25790 33182 25842 33234
rect 29262 33182 29314 33234
rect 32286 33182 32338 33234
rect 34974 33182 35026 33234
rect 35870 33182 35922 33234
rect 36206 33182 36258 33234
rect 10894 33070 10946 33122
rect 16830 33070 16882 33122
rect 18958 33070 19010 33122
rect 22430 33070 22482 33122
rect 31166 33070 31218 33122
rect 31278 33070 31330 33122
rect 31390 33070 31442 33122
rect 31614 33070 31666 33122
rect 32174 33070 32226 33122
rect 35646 33070 35698 33122
rect 35758 33070 35810 33122
rect 36318 33070 36370 33122
rect 36542 33070 36594 33122
rect 37102 33070 37154 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 8542 32734 8594 32786
rect 8766 32734 8818 32786
rect 23998 32734 24050 32786
rect 25678 32734 25730 32786
rect 26014 32734 26066 32786
rect 26910 32734 26962 32786
rect 27358 32734 27410 32786
rect 29934 32734 29986 32786
rect 33294 32734 33346 32786
rect 37102 32734 37154 32786
rect 7646 32622 7698 32674
rect 8318 32622 8370 32674
rect 10558 32622 10610 32674
rect 17726 32622 17778 32674
rect 19070 32622 19122 32674
rect 19630 32622 19682 32674
rect 24334 32622 24386 32674
rect 24558 32622 24610 32674
rect 28926 32622 28978 32674
rect 29486 32622 29538 32674
rect 31838 32622 31890 32674
rect 33630 32622 33682 32674
rect 37774 32622 37826 32674
rect 7982 32510 8034 32562
rect 8990 32510 9042 32562
rect 9662 32510 9714 32562
rect 10110 32510 10162 32562
rect 16494 32510 16546 32562
rect 17390 32510 17442 32562
rect 18622 32510 18674 32562
rect 18846 32510 18898 32562
rect 19406 32510 19458 32562
rect 19966 32510 20018 32562
rect 20526 32510 20578 32562
rect 20750 32510 20802 32562
rect 25566 32510 25618 32562
rect 25790 32510 25842 32562
rect 29038 32510 29090 32562
rect 29262 32510 29314 32562
rect 29822 32510 29874 32562
rect 30046 32510 30098 32562
rect 30494 32510 30546 32562
rect 31054 32510 31106 32562
rect 31390 32510 31442 32562
rect 34414 32510 34466 32562
rect 35982 32510 36034 32562
rect 36654 32510 36706 32562
rect 36878 32510 36930 32562
rect 37326 32510 37378 32562
rect 37662 32510 37714 32562
rect 8654 32398 8706 32450
rect 12238 32398 12290 32450
rect 19854 32398 19906 32450
rect 24670 32398 24722 32450
rect 31502 32398 31554 32450
rect 33966 32398 34018 32450
rect 34750 32398 34802 32450
rect 35310 32398 35362 32450
rect 35646 32398 35698 32450
rect 36990 32398 37042 32450
rect 19182 32286 19234 32338
rect 20638 32286 20690 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 12798 31838 12850 31890
rect 15822 31838 15874 31890
rect 18734 31838 18786 31890
rect 34638 31838 34690 31890
rect 37886 31838 37938 31890
rect 15710 31726 15762 31778
rect 16606 31726 16658 31778
rect 18510 31726 18562 31778
rect 19742 31726 19794 31778
rect 23214 31726 23266 31778
rect 23550 31726 23602 31778
rect 24110 31726 24162 31778
rect 24670 31726 24722 31778
rect 26574 31726 26626 31778
rect 27134 31726 27186 31778
rect 27582 31726 27634 31778
rect 28142 31726 28194 31778
rect 31390 31726 31442 31778
rect 33406 31726 33458 31778
rect 33742 31726 33794 31778
rect 34190 31726 34242 31778
rect 35758 31726 35810 31778
rect 36206 31726 36258 31778
rect 36878 31726 36930 31778
rect 37102 31726 37154 31778
rect 37214 31726 37266 31778
rect 38222 31726 38274 31778
rect 12686 31614 12738 31666
rect 19182 31614 19234 31666
rect 20302 31614 20354 31666
rect 21422 31614 21474 31666
rect 21534 31614 21586 31666
rect 23774 31614 23826 31666
rect 25342 31614 25394 31666
rect 27470 31614 27522 31666
rect 30830 31614 30882 31666
rect 33294 31614 33346 31666
rect 35310 31614 35362 31666
rect 37550 31614 37602 31666
rect 8318 31502 8370 31554
rect 9214 31502 9266 31554
rect 20078 31502 20130 31554
rect 20414 31502 20466 31554
rect 20862 31502 20914 31554
rect 21198 31502 21250 31554
rect 21870 31502 21922 31554
rect 22206 31502 22258 31554
rect 23550 31502 23602 31554
rect 25006 31502 25058 31554
rect 25902 31502 25954 31554
rect 26686 31502 26738 31554
rect 26798 31502 26850 31554
rect 29822 31502 29874 31554
rect 37998 31502 38050 31554
rect 38670 31502 38722 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 11678 31166 11730 31218
rect 19070 31166 19122 31218
rect 26462 31166 26514 31218
rect 26910 31166 26962 31218
rect 27246 31166 27298 31218
rect 35534 31166 35586 31218
rect 35870 31166 35922 31218
rect 36542 31166 36594 31218
rect 12910 31054 12962 31106
rect 25902 31054 25954 31106
rect 26238 31054 26290 31106
rect 35086 31054 35138 31106
rect 35310 31054 35362 31106
rect 37998 31054 38050 31106
rect 10110 30942 10162 30994
rect 11454 30942 11506 30994
rect 12238 30942 12290 30994
rect 15934 30942 15986 30994
rect 16382 30942 16434 30994
rect 19182 30942 19234 30994
rect 23886 30942 23938 30994
rect 24334 30942 24386 30994
rect 25566 30942 25618 30994
rect 26798 30942 26850 30994
rect 27246 30942 27298 30994
rect 35758 30942 35810 30994
rect 36318 30942 36370 30994
rect 37214 30942 37266 30994
rect 15038 30830 15090 30882
rect 16830 30830 16882 30882
rect 17502 30830 17554 30882
rect 30270 30830 30322 30882
rect 35646 30830 35698 30882
rect 40126 30830 40178 30882
rect 9550 30718 9602 30770
rect 9886 30718 9938 30770
rect 19070 30718 19122 30770
rect 26574 30718 26626 30770
rect 36654 30718 36706 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 27582 30382 27634 30434
rect 27806 30382 27858 30434
rect 37662 30382 37714 30434
rect 8206 30270 8258 30322
rect 8990 30270 9042 30322
rect 10894 30270 10946 30322
rect 22990 30270 23042 30322
rect 30718 30270 30770 30322
rect 31278 30270 31330 30322
rect 32062 30270 32114 30322
rect 32398 30270 32450 30322
rect 34638 30270 34690 30322
rect 36318 30270 36370 30322
rect 37998 30270 38050 30322
rect 8542 30158 8594 30210
rect 9550 30158 9602 30210
rect 9886 30158 9938 30210
rect 17838 30158 17890 30210
rect 17950 30158 18002 30210
rect 18174 30158 18226 30210
rect 18398 30158 18450 30210
rect 22766 30158 22818 30210
rect 23326 30158 23378 30210
rect 25902 30158 25954 30210
rect 26462 30158 26514 30210
rect 27134 30158 27186 30210
rect 28030 30158 28082 30210
rect 28366 30158 28418 30210
rect 29262 30158 29314 30210
rect 31838 30158 31890 30210
rect 32958 30158 33010 30210
rect 33966 30158 34018 30210
rect 37326 30158 37378 30210
rect 7870 30046 7922 30098
rect 9998 30046 10050 30098
rect 18734 30046 18786 30098
rect 19182 30046 19234 30098
rect 20862 30046 20914 30098
rect 22206 30046 22258 30098
rect 26238 30046 26290 30098
rect 26910 30046 26962 30098
rect 29486 30046 29538 30098
rect 30382 30046 30434 30098
rect 32174 30046 32226 30098
rect 34414 30046 34466 30098
rect 34526 30046 34578 30098
rect 36990 30046 37042 30098
rect 8094 29934 8146 29986
rect 8318 29934 8370 29986
rect 9438 29934 9490 29986
rect 12350 29934 12402 29986
rect 18510 29934 18562 29986
rect 18622 29934 18674 29986
rect 18958 29934 19010 29986
rect 21534 29934 21586 29986
rect 21870 29934 21922 29986
rect 26014 29934 26066 29986
rect 28478 29934 28530 29986
rect 28702 29934 28754 29986
rect 30606 29934 30658 29986
rect 30830 29934 30882 29986
rect 31166 29934 31218 29986
rect 31390 29934 31442 29986
rect 32622 29934 32674 29986
rect 32846 29934 32898 29986
rect 33630 29934 33682 29986
rect 35982 29934 36034 29986
rect 36430 29934 36482 29986
rect 37886 29934 37938 29986
rect 38446 29934 38498 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 16718 29598 16770 29650
rect 18958 29598 19010 29650
rect 29598 29598 29650 29650
rect 31950 29598 32002 29650
rect 36094 29598 36146 29650
rect 7982 29486 8034 29538
rect 17502 29486 17554 29538
rect 19294 29486 19346 29538
rect 20750 29486 20802 29538
rect 21198 29486 21250 29538
rect 26574 29486 26626 29538
rect 26910 29486 26962 29538
rect 27022 29486 27074 29538
rect 29486 29486 29538 29538
rect 30606 29486 30658 29538
rect 31838 29486 31890 29538
rect 37998 29486 38050 29538
rect 8654 29374 8706 29426
rect 8878 29374 8930 29426
rect 9662 29374 9714 29426
rect 9774 29374 9826 29426
rect 10222 29374 10274 29426
rect 13582 29374 13634 29426
rect 16830 29374 16882 29426
rect 17390 29374 17442 29426
rect 18286 29374 18338 29426
rect 18510 29374 18562 29426
rect 19182 29374 19234 29426
rect 20862 29374 20914 29426
rect 21422 29374 21474 29426
rect 21758 29374 21810 29426
rect 22766 29374 22818 29426
rect 23326 29374 23378 29426
rect 24110 29374 24162 29426
rect 26686 29374 26738 29426
rect 30830 29374 30882 29426
rect 33070 29374 33122 29426
rect 33294 29374 33346 29426
rect 35534 29374 35586 29426
rect 35870 29374 35922 29426
rect 37214 29374 37266 29426
rect 9998 29262 10050 29314
rect 10782 29262 10834 29314
rect 12910 29262 12962 29314
rect 14478 29262 14530 29314
rect 18062 29262 18114 29314
rect 20078 29262 20130 29314
rect 23774 29262 23826 29314
rect 33854 29262 33906 29314
rect 35982 29262 36034 29314
rect 36878 29262 36930 29314
rect 40126 29262 40178 29314
rect 16718 29150 16770 29202
rect 17502 29150 17554 29202
rect 29598 29150 29650 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 5966 28814 6018 28866
rect 19630 28814 19682 28866
rect 19854 28814 19906 28866
rect 5630 28702 5682 28754
rect 7086 28702 7138 28754
rect 9214 28702 9266 28754
rect 9550 28702 9602 28754
rect 10446 28702 10498 28754
rect 11118 28702 11170 28754
rect 15374 28702 15426 28754
rect 17054 28702 17106 28754
rect 18062 28702 18114 28754
rect 24222 28702 24274 28754
rect 25902 28702 25954 28754
rect 28030 28702 28082 28754
rect 28478 28702 28530 28754
rect 31502 28702 31554 28754
rect 6302 28590 6354 28642
rect 10222 28590 10274 28642
rect 11566 28590 11618 28642
rect 12574 28590 12626 28642
rect 13806 28590 13858 28642
rect 13918 28590 13970 28642
rect 14814 28590 14866 28642
rect 15710 28590 15762 28642
rect 16830 28590 16882 28642
rect 18174 28590 18226 28642
rect 18734 28590 18786 28642
rect 19406 28590 19458 28642
rect 23662 28590 23714 28642
rect 24894 28590 24946 28642
rect 25230 28590 25282 28642
rect 31278 28590 31330 28642
rect 35422 28590 35474 28642
rect 38558 28590 38610 28642
rect 12014 28478 12066 28530
rect 13470 28478 13522 28530
rect 14142 28478 14194 28530
rect 14254 28478 14306 28530
rect 17726 28478 17778 28530
rect 31726 28478 31778 28530
rect 38222 28478 38274 28530
rect 5742 28366 5794 28418
rect 12350 28366 12402 28418
rect 13582 28366 13634 28418
rect 19518 28366 19570 28418
rect 22430 28366 22482 28418
rect 24110 28366 24162 28418
rect 24334 28366 24386 28418
rect 35534 28366 35586 28418
rect 35758 28366 35810 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 9662 28030 9714 28082
rect 18398 28030 18450 28082
rect 33070 28030 33122 28082
rect 5406 27918 5458 27970
rect 17838 27918 17890 27970
rect 18510 27918 18562 27970
rect 22542 27918 22594 27970
rect 27358 27918 27410 27970
rect 27918 27918 27970 27970
rect 32286 27918 32338 27970
rect 4734 27806 4786 27858
rect 9550 27806 9602 27858
rect 9774 27806 9826 27858
rect 10222 27806 10274 27858
rect 15934 27806 15986 27858
rect 16382 27806 16434 27858
rect 17502 27806 17554 27858
rect 18174 27806 18226 27858
rect 18846 27806 18898 27858
rect 22878 27806 22930 27858
rect 27582 27806 27634 27858
rect 28254 27806 28306 27858
rect 31838 27806 31890 27858
rect 32062 27806 32114 27858
rect 33294 27806 33346 27858
rect 33518 27806 33570 27858
rect 35870 27806 35922 27858
rect 7534 27694 7586 27746
rect 13358 27694 13410 27746
rect 17614 27694 17666 27746
rect 18958 27694 19010 27746
rect 19406 27694 19458 27746
rect 25342 27694 25394 27746
rect 35422 27694 35474 27746
rect 36318 27694 36370 27746
rect 27246 27582 27298 27634
rect 31950 27582 32002 27634
rect 32958 27582 33010 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 10334 27246 10386 27298
rect 11006 27246 11058 27298
rect 17166 27246 17218 27298
rect 31950 27246 32002 27298
rect 32174 27246 32226 27298
rect 33854 27246 33906 27298
rect 35310 27246 35362 27298
rect 37998 27246 38050 27298
rect 6974 27134 7026 27186
rect 10558 27134 10610 27186
rect 11006 27134 11058 27186
rect 12126 27134 12178 27186
rect 12910 27134 12962 27186
rect 15934 27134 15986 27186
rect 18286 27134 18338 27186
rect 21310 27134 21362 27186
rect 24670 27134 24722 27186
rect 25790 27134 25842 27186
rect 26686 27134 26738 27186
rect 27694 27134 27746 27186
rect 28030 27134 28082 27186
rect 29822 27134 29874 27186
rect 31614 27134 31666 27186
rect 32958 27134 33010 27186
rect 34862 27134 34914 27186
rect 38558 27134 38610 27186
rect 6526 27022 6578 27074
rect 12462 27022 12514 27074
rect 16158 27022 16210 27074
rect 16830 27022 16882 27074
rect 17502 27022 17554 27074
rect 19294 27022 19346 27074
rect 19518 27022 19570 27074
rect 19742 27022 19794 27074
rect 20190 27022 20242 27074
rect 20414 27022 20466 27074
rect 20638 27022 20690 27074
rect 24222 27022 24274 27074
rect 26238 27022 26290 27074
rect 27582 27022 27634 27074
rect 29038 27022 29090 27074
rect 29486 27022 29538 27074
rect 29598 27022 29650 27074
rect 30046 27022 30098 27074
rect 31502 27022 31554 27074
rect 32846 27022 32898 27074
rect 33294 27022 33346 27074
rect 34302 27022 34354 27074
rect 35422 27022 35474 27074
rect 35982 27022 36034 27074
rect 38334 27022 38386 27074
rect 39566 27022 39618 27074
rect 40014 27022 40066 27074
rect 6190 26910 6242 26962
rect 18398 26910 18450 26962
rect 18622 26910 18674 26962
rect 20750 26910 20802 26962
rect 23438 26910 23490 26962
rect 28590 26910 28642 26962
rect 31390 26910 31442 26962
rect 33070 26910 33122 26962
rect 34526 26910 34578 26962
rect 34750 26910 34802 26962
rect 17614 26798 17666 26850
rect 17726 26798 17778 26850
rect 17838 26798 17890 26850
rect 19630 26798 19682 26850
rect 29486 26798 29538 26850
rect 32734 26798 32786 26850
rect 39790 26798 39842 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 19182 26462 19234 26514
rect 19966 26462 20018 26514
rect 23550 26462 23602 26514
rect 31390 26462 31442 26514
rect 33294 26462 33346 26514
rect 39566 26462 39618 26514
rect 2046 26350 2098 26402
rect 3950 26350 4002 26402
rect 19294 26350 19346 26402
rect 28366 26350 28418 26402
rect 33070 26350 33122 26402
rect 34862 26350 34914 26402
rect 36318 26350 36370 26402
rect 39790 26350 39842 26402
rect 40126 26350 40178 26402
rect 1822 26238 1874 26290
rect 23214 26238 23266 26290
rect 24334 26238 24386 26290
rect 27694 26238 27746 26290
rect 30942 26238 30994 26290
rect 31726 26238 31778 26290
rect 32062 26238 32114 26290
rect 32286 26238 32338 26290
rect 33294 26238 33346 26290
rect 33854 26238 33906 26290
rect 35758 26238 35810 26290
rect 36430 26238 36482 26290
rect 36766 26238 36818 26290
rect 2494 26126 2546 26178
rect 20974 26126 21026 26178
rect 24558 26126 24610 26178
rect 26910 26126 26962 26178
rect 30494 26126 30546 26178
rect 35310 26126 35362 26178
rect 3838 26014 3890 26066
rect 4174 26014 4226 26066
rect 23998 26014 24050 26066
rect 30718 26014 30770 26066
rect 31278 26014 31330 26066
rect 31502 26014 31554 26066
rect 33518 26014 33570 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 24334 25678 24386 25730
rect 1710 25566 1762 25618
rect 3838 25566 3890 25618
rect 10334 25566 10386 25618
rect 11454 25566 11506 25618
rect 16382 25566 16434 25618
rect 23886 25566 23938 25618
rect 31166 25566 31218 25618
rect 32174 25566 32226 25618
rect 32958 25566 33010 25618
rect 34078 25566 34130 25618
rect 34750 25566 34802 25618
rect 35646 25566 35698 25618
rect 4622 25454 4674 25506
rect 10110 25454 10162 25506
rect 13470 25454 13522 25506
rect 18846 25454 18898 25506
rect 24782 25454 24834 25506
rect 30270 25454 30322 25506
rect 31054 25454 31106 25506
rect 32510 25454 32562 25506
rect 33742 25454 33794 25506
rect 35198 25454 35250 25506
rect 10222 25342 10274 25394
rect 10894 25342 10946 25394
rect 14254 25342 14306 25394
rect 19182 25342 19234 25394
rect 22766 25342 22818 25394
rect 23774 25342 23826 25394
rect 24222 25342 24274 25394
rect 29486 25342 29538 25394
rect 29710 25342 29762 25394
rect 29934 25342 29986 25394
rect 31614 25342 31666 25394
rect 33294 25342 33346 25394
rect 9214 25230 9266 25282
rect 11006 25230 11058 25282
rect 22430 25230 22482 25282
rect 25006 25230 25058 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 6526 24894 6578 24946
rect 10782 24894 10834 24946
rect 31838 24894 31890 24946
rect 33406 24894 33458 24946
rect 33518 24894 33570 24946
rect 33630 24894 33682 24946
rect 36878 24894 36930 24946
rect 5294 24782 5346 24834
rect 6862 24782 6914 24834
rect 22318 24782 22370 24834
rect 30830 24782 30882 24834
rect 32286 24782 32338 24834
rect 4622 24670 4674 24722
rect 5070 24670 5122 24722
rect 6302 24670 6354 24722
rect 6414 24670 6466 24722
rect 6638 24670 6690 24722
rect 7310 24670 7362 24722
rect 7422 24670 7474 24722
rect 7646 24670 7698 24722
rect 7758 24670 7810 24722
rect 8654 24670 8706 24722
rect 9774 24670 9826 24722
rect 10334 24670 10386 24722
rect 10670 24670 10722 24722
rect 11566 24670 11618 24722
rect 17502 24670 17554 24722
rect 17838 24670 17890 24722
rect 18062 24670 18114 24722
rect 21198 24670 21250 24722
rect 22094 24670 22146 24722
rect 25790 24670 25842 24722
rect 26126 24670 26178 24722
rect 26686 24670 26738 24722
rect 31390 24670 31442 24722
rect 32398 24670 32450 24722
rect 32958 24670 33010 24722
rect 37214 24670 37266 24722
rect 1710 24558 1762 24610
rect 3838 24558 3890 24610
rect 7534 24558 7586 24610
rect 12350 24558 12402 24610
rect 14478 24558 14530 24610
rect 17614 24558 17666 24610
rect 20862 24558 20914 24610
rect 25230 24558 25282 24610
rect 37998 24558 38050 24610
rect 40126 24558 40178 24610
rect 8654 24446 8706 24498
rect 8990 24446 9042 24498
rect 10782 24446 10834 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3838 24110 3890 24162
rect 4174 24110 4226 24162
rect 23886 24110 23938 24162
rect 1934 23998 1986 24050
rect 8542 23998 8594 24050
rect 10670 23998 10722 24050
rect 18062 23998 18114 24050
rect 18958 23998 19010 24050
rect 20190 23998 20242 24050
rect 20750 23998 20802 24050
rect 40126 23998 40178 24050
rect 2942 23886 2994 23938
rect 3838 23886 3890 23938
rect 6750 23886 6802 23938
rect 7982 23886 8034 23938
rect 11454 23886 11506 23938
rect 16606 23886 16658 23938
rect 17054 23886 17106 23938
rect 17278 23886 17330 23938
rect 17726 23886 17778 23938
rect 18510 23886 18562 23938
rect 19854 23886 19906 23938
rect 22318 23886 22370 23938
rect 23102 23886 23154 23938
rect 23662 23886 23714 23938
rect 24222 23886 24274 23938
rect 36542 23886 36594 23938
rect 37214 23886 37266 23938
rect 6414 23774 6466 23826
rect 19630 23774 19682 23826
rect 20190 23774 20242 23826
rect 20638 23774 20690 23826
rect 22766 23774 22818 23826
rect 24446 23774 24498 23826
rect 37998 23774 38050 23826
rect 6526 23662 6578 23714
rect 7758 23662 7810 23714
rect 16382 23662 16434 23714
rect 17502 23662 17554 23714
rect 17950 23662 18002 23714
rect 18174 23662 18226 23714
rect 20078 23662 20130 23714
rect 21870 23662 21922 23714
rect 22094 23662 22146 23714
rect 22878 23662 22930 23714
rect 24334 23662 24386 23714
rect 29822 23662 29874 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 4734 23326 4786 23378
rect 5294 23326 5346 23378
rect 6526 23326 6578 23378
rect 7198 23326 7250 23378
rect 36654 23326 36706 23378
rect 37550 23326 37602 23378
rect 4510 23214 4562 23266
rect 5070 23214 5122 23266
rect 5966 23214 6018 23266
rect 7422 23214 7474 23266
rect 8878 23214 8930 23266
rect 15486 23214 15538 23266
rect 16382 23214 16434 23266
rect 18062 23214 18114 23266
rect 23326 23214 23378 23266
rect 30046 23214 30098 23266
rect 34414 23214 34466 23266
rect 36318 23214 36370 23266
rect 37438 23214 37490 23266
rect 4398 23102 4450 23154
rect 4958 23102 5010 23154
rect 5518 23102 5570 23154
rect 5630 23102 5682 23154
rect 5742 23102 5794 23154
rect 7086 23102 7138 23154
rect 10334 23102 10386 23154
rect 12350 23102 12402 23154
rect 13022 23102 13074 23154
rect 15822 23102 15874 23154
rect 16270 23102 16322 23154
rect 17726 23102 17778 23154
rect 17950 23102 18002 23154
rect 18510 23102 18562 23154
rect 19518 23102 19570 23154
rect 26574 23102 26626 23154
rect 29822 23102 29874 23154
rect 30494 23102 30546 23154
rect 34302 23102 34354 23154
rect 34638 23102 34690 23154
rect 9886 22990 9938 23042
rect 15150 22990 15202 23042
rect 16158 22990 16210 23042
rect 19070 22990 19122 23042
rect 27358 22990 27410 23042
rect 29486 22990 29538 23042
rect 29934 22990 29986 23042
rect 6414 22878 6466 22930
rect 6750 22878 6802 22930
rect 8654 22878 8706 22930
rect 8990 22878 9042 22930
rect 17614 22878 17666 22930
rect 18510 22878 18562 22930
rect 18958 22878 19010 22930
rect 37662 22878 37714 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 16494 22542 16546 22594
rect 29038 22542 29090 22594
rect 33742 22542 33794 22594
rect 5070 22430 5122 22482
rect 6414 22430 6466 22482
rect 11342 22430 11394 22482
rect 12126 22430 12178 22482
rect 15710 22430 15762 22482
rect 22990 22430 23042 22482
rect 25118 22430 25170 22482
rect 27358 22430 27410 22482
rect 28142 22430 28194 22482
rect 33406 22430 33458 22482
rect 4734 22318 4786 22370
rect 6302 22318 6354 22370
rect 11678 22318 11730 22370
rect 15374 22318 15426 22370
rect 15934 22318 15986 22370
rect 16270 22318 16322 22370
rect 16718 22318 16770 22370
rect 19630 22318 19682 22370
rect 21646 22318 21698 22370
rect 25790 22318 25842 22370
rect 26350 22318 26402 22370
rect 26798 22318 26850 22370
rect 27470 22318 27522 22370
rect 27806 22318 27858 22370
rect 28254 22318 28306 22370
rect 29374 22318 29426 22370
rect 35310 22318 35362 22370
rect 35870 22318 35922 22370
rect 37326 22318 37378 22370
rect 37886 22318 37938 22370
rect 38222 22318 38274 22370
rect 4958 22206 5010 22258
rect 6190 22206 6242 22258
rect 18286 22206 18338 22258
rect 21310 22206 21362 22258
rect 28030 22206 28082 22258
rect 28478 22206 28530 22258
rect 29598 22206 29650 22258
rect 32734 22206 32786 22258
rect 33070 22206 33122 22258
rect 34190 22206 34242 22258
rect 34414 22206 34466 22258
rect 35534 22206 35586 22258
rect 36206 22206 36258 22258
rect 37998 22206 38050 22258
rect 38558 22206 38610 22258
rect 6526 22094 6578 22146
rect 6750 22094 6802 22146
rect 17166 22094 17218 22146
rect 17950 22094 18002 22146
rect 19294 22094 19346 22146
rect 27246 22094 27298 22146
rect 29150 22094 29202 22146
rect 33518 22094 33570 22146
rect 34526 22094 34578 22146
rect 34638 22094 34690 22146
rect 36094 22094 36146 22146
rect 38446 22094 38498 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 3054 21758 3106 21810
rect 3502 21758 3554 21810
rect 4846 21758 4898 21810
rect 5406 21758 5458 21810
rect 6750 21758 6802 21810
rect 6862 21758 6914 21810
rect 7198 21758 7250 21810
rect 26910 21758 26962 21810
rect 28926 21758 28978 21810
rect 36430 21758 36482 21810
rect 37886 21758 37938 21810
rect 2942 21646 2994 21698
rect 3838 21646 3890 21698
rect 6638 21646 6690 21698
rect 7534 21646 7586 21698
rect 13918 21646 13970 21698
rect 15374 21646 15426 21698
rect 15710 21646 15762 21698
rect 16382 21646 16434 21698
rect 19294 21646 19346 21698
rect 27918 21646 27970 21698
rect 28142 21646 28194 21698
rect 29598 21646 29650 21698
rect 32174 21646 32226 21698
rect 33070 21646 33122 21698
rect 33406 21646 33458 21698
rect 34862 21646 34914 21698
rect 35198 21646 35250 21698
rect 37550 21646 37602 21698
rect 4622 21534 4674 21586
rect 5182 21534 5234 21586
rect 5630 21534 5682 21586
rect 5966 21534 6018 21586
rect 6190 21534 6242 21586
rect 13582 21534 13634 21586
rect 15262 21534 15314 21586
rect 16158 21534 16210 21586
rect 16270 21534 16322 21586
rect 18174 21534 18226 21586
rect 23774 21534 23826 21586
rect 27582 21534 27634 21586
rect 28814 21534 28866 21586
rect 29486 21534 29538 21586
rect 31502 21534 31554 21586
rect 32510 21534 32562 21586
rect 33182 21534 33234 21586
rect 33630 21534 33682 21586
rect 35422 21534 35474 21586
rect 35870 21534 35922 21586
rect 36990 21534 37042 21586
rect 37214 21534 37266 21586
rect 38110 21534 38162 21586
rect 39118 21534 39170 21586
rect 5518 21422 5570 21474
rect 15598 21422 15650 21474
rect 16830 21422 16882 21474
rect 17950 21422 18002 21474
rect 19406 21422 19458 21474
rect 20862 21422 20914 21474
rect 22990 21422 23042 21474
rect 24222 21422 24274 21474
rect 26126 21422 26178 21474
rect 27694 21422 27746 21474
rect 30158 21422 30210 21474
rect 34190 21422 34242 21474
rect 40014 21422 40066 21474
rect 3054 21310 3106 21362
rect 18398 21310 18450 21362
rect 18846 21310 18898 21362
rect 19070 21310 19122 21362
rect 29598 21310 29650 21362
rect 31502 21310 31554 21362
rect 31838 21310 31890 21362
rect 33854 21310 33906 21362
rect 36094 21310 36146 21362
rect 37438 21310 37490 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 4958 20974 5010 21026
rect 5742 20974 5794 21026
rect 5854 20974 5906 21026
rect 16718 20974 16770 21026
rect 21534 20974 21586 21026
rect 21870 20974 21922 21026
rect 30830 20974 30882 21026
rect 6862 20862 6914 20914
rect 11678 20862 11730 20914
rect 12014 20862 12066 20914
rect 18846 20862 18898 20914
rect 40126 20862 40178 20914
rect 3614 20750 3666 20802
rect 6078 20750 6130 20802
rect 6190 20750 6242 20802
rect 6638 20750 6690 20802
rect 10110 20750 10162 20802
rect 12238 20750 12290 20802
rect 17278 20750 17330 20802
rect 17838 20750 17890 20802
rect 18062 20750 18114 20802
rect 20078 20750 20130 20802
rect 21310 20750 21362 20802
rect 21758 20750 21810 20802
rect 29486 20750 29538 20802
rect 29710 20750 29762 20802
rect 31278 20750 31330 20802
rect 31502 20750 31554 20802
rect 31614 20750 31666 20802
rect 31726 20750 31778 20802
rect 32174 20750 32226 20802
rect 34190 20750 34242 20802
rect 37214 20750 37266 20802
rect 1710 20638 1762 20690
rect 3166 20638 3218 20690
rect 5070 20638 5122 20690
rect 6974 20638 7026 20690
rect 9214 20638 9266 20690
rect 9550 20638 9602 20690
rect 11342 20638 11394 20690
rect 11566 20638 11618 20690
rect 13470 20638 13522 20690
rect 13582 20638 13634 20690
rect 16046 20638 16098 20690
rect 16382 20638 16434 20690
rect 17166 20638 17218 20690
rect 17390 20638 17442 20690
rect 18174 20638 18226 20690
rect 19518 20638 19570 20690
rect 19742 20638 19794 20690
rect 29150 20638 29202 20690
rect 33294 20638 33346 20690
rect 34750 20638 34802 20690
rect 37998 20638 38050 20690
rect 2046 20526 2098 20578
rect 2494 20526 2546 20578
rect 2942 20526 2994 20578
rect 3054 20526 3106 20578
rect 3838 20526 3890 20578
rect 4174 20526 4226 20578
rect 4510 20526 4562 20578
rect 4958 20526 5010 20578
rect 9886 20526 9938 20578
rect 12574 20526 12626 20578
rect 13806 20526 13858 20578
rect 18622 20526 18674 20578
rect 29262 20526 29314 20578
rect 33630 20526 33682 20578
rect 36430 20526 36482 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 2382 20190 2434 20242
rect 3838 20190 3890 20242
rect 5630 20190 5682 20242
rect 5742 20190 5794 20242
rect 6862 20190 6914 20242
rect 8430 20190 8482 20242
rect 17950 20190 18002 20242
rect 18174 20190 18226 20242
rect 20974 20190 21026 20242
rect 25790 20190 25842 20242
rect 33406 20190 33458 20242
rect 34750 20190 34802 20242
rect 3278 20078 3330 20130
rect 3726 20078 3778 20130
rect 5294 20078 5346 20130
rect 6638 20078 6690 20130
rect 11790 20078 11842 20130
rect 12014 20078 12066 20130
rect 13134 20078 13186 20130
rect 13358 20078 13410 20130
rect 13918 20078 13970 20130
rect 14478 20078 14530 20130
rect 14590 20078 14642 20130
rect 19294 20078 19346 20130
rect 20414 20078 20466 20130
rect 21646 20078 21698 20130
rect 26126 20078 26178 20130
rect 27582 20078 27634 20130
rect 34302 20078 34354 20130
rect 2158 19966 2210 20018
rect 2718 19966 2770 20018
rect 4286 19966 4338 20018
rect 4734 19966 4786 20018
rect 5854 19966 5906 20018
rect 6190 19966 6242 20018
rect 6526 19966 6578 20018
rect 8206 19966 8258 20018
rect 8542 19966 8594 20018
rect 8654 19966 8706 20018
rect 8990 19966 9042 20018
rect 10334 19966 10386 20018
rect 12238 19966 12290 20018
rect 12574 19966 12626 20018
rect 12798 19966 12850 20018
rect 13470 19966 13522 20018
rect 13694 19966 13746 20018
rect 14254 19966 14306 20018
rect 17838 19966 17890 20018
rect 19630 19966 19682 20018
rect 20190 19966 20242 20018
rect 20638 19966 20690 20018
rect 20750 19966 20802 20018
rect 21198 19966 21250 20018
rect 21870 19966 21922 20018
rect 26350 19966 26402 20018
rect 26686 19966 26738 20018
rect 27246 19966 27298 20018
rect 29934 19966 29986 20018
rect 31838 19966 31890 20018
rect 32062 19966 32114 20018
rect 32510 19966 32562 20018
rect 33518 19966 33570 20018
rect 33742 19966 33794 20018
rect 34078 19966 34130 20018
rect 34638 20022 34690 20074
rect 38894 20078 38946 20130
rect 39678 20078 39730 20130
rect 34862 19966 34914 20018
rect 35086 19966 35138 20018
rect 35422 19966 35474 20018
rect 37102 19966 37154 20018
rect 9662 19854 9714 19906
rect 10110 19854 10162 19906
rect 11006 19854 11058 19906
rect 12014 19854 12066 19906
rect 18958 19854 19010 19906
rect 21422 19854 21474 19906
rect 25230 19854 25282 19906
rect 26462 19854 26514 19906
rect 27470 19854 27522 19906
rect 31278 19854 31330 19906
rect 37326 19854 37378 19906
rect 14030 19742 14082 19794
rect 32286 19742 32338 19794
rect 37886 19742 37938 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 3278 19406 3330 19458
rect 5742 19406 5794 19458
rect 10782 19406 10834 19458
rect 11118 19406 11170 19458
rect 12014 19406 12066 19458
rect 12798 19406 12850 19458
rect 15038 19406 15090 19458
rect 20750 19406 20802 19458
rect 21422 19406 21474 19458
rect 23774 19406 23826 19458
rect 37774 19406 37826 19458
rect 2494 19294 2546 19346
rect 3054 19294 3106 19346
rect 4734 19294 4786 19346
rect 9550 19294 9602 19346
rect 10558 19294 10610 19346
rect 13582 19294 13634 19346
rect 14478 19294 14530 19346
rect 21758 19294 21810 19346
rect 28142 19294 28194 19346
rect 37998 19294 38050 19346
rect 40014 19294 40066 19346
rect 1710 19182 1762 19234
rect 4174 19182 4226 19234
rect 4622 19182 4674 19234
rect 5630 19182 5682 19234
rect 7870 19182 7922 19234
rect 8318 19182 8370 19234
rect 8990 19182 9042 19234
rect 9438 19182 9490 19234
rect 12574 19182 12626 19234
rect 14030 19182 14082 19234
rect 14814 19182 14866 19234
rect 15374 19182 15426 19234
rect 18510 19182 18562 19234
rect 18958 19182 19010 19234
rect 19966 19182 20018 19234
rect 24334 19182 24386 19234
rect 24670 19182 24722 19234
rect 25230 19182 25282 19234
rect 28590 19182 28642 19234
rect 30382 19182 30434 19234
rect 32622 19182 32674 19234
rect 37438 19182 37490 19234
rect 38894 19182 38946 19234
rect 2046 19070 2098 19122
rect 6302 19070 6354 19122
rect 7310 19070 7362 19122
rect 7534 19070 7586 19122
rect 9662 19070 9714 19122
rect 12238 19070 12290 19122
rect 17278 19070 17330 19122
rect 17614 19070 17666 19122
rect 18062 19070 18114 19122
rect 19518 19070 19570 19122
rect 20190 19070 20242 19122
rect 20302 19070 20354 19122
rect 21646 19070 21698 19122
rect 23886 19070 23938 19122
rect 24894 19070 24946 19122
rect 26014 19070 26066 19122
rect 29486 19070 29538 19122
rect 30606 19070 30658 19122
rect 31278 19070 31330 19122
rect 31614 19070 31666 19122
rect 32958 19070 33010 19122
rect 3614 18958 3666 19010
rect 6414 18958 6466 19010
rect 6638 18958 6690 19010
rect 7758 18958 7810 19010
rect 8206 18958 8258 19010
rect 8430 18958 8482 19010
rect 8654 18958 8706 19010
rect 12910 18958 12962 19010
rect 19406 18958 19458 19010
rect 24782 18958 24834 19010
rect 29822 18958 29874 19010
rect 30942 18958 30994 19010
rect 31950 18958 32002 19010
rect 37102 18958 37154 19010
rect 37998 18958 38050 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 3838 18622 3890 18674
rect 4286 18622 4338 18674
rect 5182 18622 5234 18674
rect 5294 18622 5346 18674
rect 7422 18622 7474 18674
rect 8206 18622 8258 18674
rect 8990 18622 9042 18674
rect 13918 18622 13970 18674
rect 18846 18622 18898 18674
rect 20078 18622 20130 18674
rect 20974 18622 21026 18674
rect 33742 18622 33794 18674
rect 37326 18622 37378 18674
rect 6078 18510 6130 18562
rect 6302 18510 6354 18562
rect 7646 18510 7698 18562
rect 12910 18510 12962 18562
rect 13246 18510 13298 18562
rect 14142 18510 14194 18562
rect 19742 18510 19794 18562
rect 25566 18510 25618 18562
rect 26350 18510 26402 18562
rect 29262 18510 29314 18562
rect 34638 18510 34690 18562
rect 36654 18510 36706 18562
rect 3726 18398 3778 18450
rect 4174 18398 4226 18450
rect 4510 18398 4562 18450
rect 5518 18398 5570 18450
rect 5854 18398 5906 18450
rect 7198 18398 7250 18450
rect 7870 18398 7922 18450
rect 8206 18398 8258 18450
rect 8430 18398 8482 18450
rect 13694 18398 13746 18450
rect 17838 18398 17890 18450
rect 18286 18398 18338 18450
rect 21534 18398 21586 18450
rect 22206 18398 22258 18450
rect 25342 18398 25394 18450
rect 26574 18398 26626 18450
rect 27246 18398 27298 18450
rect 34078 18398 34130 18450
rect 34414 18398 34466 18450
rect 35086 18398 35138 18450
rect 36094 18398 36146 18450
rect 36542 18398 36594 18450
rect 38894 18398 38946 18450
rect 39678 18398 39730 18450
rect 7310 18286 7362 18338
rect 24334 18286 24386 18338
rect 25678 18286 25730 18338
rect 34862 18286 34914 18338
rect 35310 18286 35362 18338
rect 35534 18286 35586 18338
rect 36318 18286 36370 18338
rect 6414 18174 6466 18226
rect 14254 18174 14306 18226
rect 18398 18174 18450 18226
rect 18846 18174 18898 18226
rect 26910 18174 26962 18226
rect 38110 18174 38162 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 17166 17838 17218 17890
rect 17838 17838 17890 17890
rect 19070 17838 19122 17890
rect 34526 17838 34578 17890
rect 19518 17726 19570 17778
rect 24558 17726 24610 17778
rect 25006 17726 25058 17778
rect 27022 17726 27074 17778
rect 27470 17726 27522 17778
rect 35534 17726 35586 17778
rect 37774 17726 37826 17778
rect 5966 17614 6018 17666
rect 6862 17614 6914 17666
rect 7198 17614 7250 17666
rect 16830 17614 16882 17666
rect 17166 17614 17218 17666
rect 18398 17614 18450 17666
rect 18622 17614 18674 17666
rect 19742 17614 19794 17666
rect 20078 17614 20130 17666
rect 27694 17614 27746 17666
rect 28254 17614 28306 17666
rect 29150 17614 29202 17666
rect 30718 17614 30770 17666
rect 31838 17614 31890 17666
rect 32398 17614 32450 17666
rect 33966 17614 34018 17666
rect 35646 17614 35698 17666
rect 37102 17614 37154 17666
rect 6190 17502 6242 17554
rect 6974 17502 7026 17554
rect 16606 17502 16658 17554
rect 18286 17502 18338 17554
rect 18958 17502 19010 17554
rect 19518 17502 19570 17554
rect 27134 17502 27186 17554
rect 27918 17502 27970 17554
rect 30158 17502 30210 17554
rect 30494 17502 30546 17554
rect 31166 17502 31218 17554
rect 31502 17502 31554 17554
rect 32622 17502 32674 17554
rect 32734 17502 32786 17554
rect 33854 17502 33906 17554
rect 34078 17502 34130 17554
rect 36318 17502 36370 17554
rect 16718 17390 16770 17442
rect 26686 17390 26738 17442
rect 28478 17390 28530 17442
rect 29486 17390 29538 17442
rect 29822 17390 29874 17442
rect 32174 17390 32226 17442
rect 40014 17390 40066 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4398 17054 4450 17106
rect 6526 17054 6578 17106
rect 16494 17054 16546 17106
rect 33406 17054 33458 17106
rect 34078 17054 34130 17106
rect 36766 17054 36818 17106
rect 4734 16942 4786 16994
rect 5742 16942 5794 16994
rect 6302 16942 6354 16994
rect 15486 16942 15538 16994
rect 16718 16942 16770 16994
rect 17726 16942 17778 16994
rect 29150 16942 29202 16994
rect 29486 16942 29538 16994
rect 30158 16942 30210 16994
rect 30494 16942 30546 16994
rect 30830 16942 30882 16994
rect 33070 16942 33122 16994
rect 36542 16942 36594 16994
rect 36654 16942 36706 16994
rect 37998 16942 38050 16994
rect 3278 16830 3330 16882
rect 5630 16830 5682 16882
rect 5966 16830 6018 16882
rect 6190 16830 6242 16882
rect 7310 16830 7362 16882
rect 7534 16830 7586 16882
rect 7758 16830 7810 16882
rect 8206 16830 8258 16882
rect 8766 16830 8818 16882
rect 16270 16830 16322 16882
rect 16830 16830 16882 16882
rect 19630 16830 19682 16882
rect 29934 16830 29986 16882
rect 34638 16830 34690 16882
rect 34974 16830 35026 16882
rect 35534 16830 35586 16882
rect 37214 16830 37266 16882
rect 7646 16718 7698 16770
rect 13358 16718 13410 16770
rect 17950 16718 18002 16770
rect 19294 16718 19346 16770
rect 34414 16718 34466 16770
rect 35198 16718 35250 16770
rect 36206 16718 36258 16770
rect 40126 16718 40178 16770
rect 3278 16606 3330 16658
rect 3614 16606 3666 16658
rect 7086 16606 7138 16658
rect 8430 16606 8482 16658
rect 18174 16606 18226 16658
rect 18398 16606 18450 16658
rect 18846 16606 18898 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 5518 16270 5570 16322
rect 6190 16270 6242 16322
rect 6750 16270 6802 16322
rect 7086 16270 7138 16322
rect 16942 16270 16994 16322
rect 17614 16270 17666 16322
rect 17950 16270 18002 16322
rect 33518 16270 33570 16322
rect 33854 16270 33906 16322
rect 34638 16270 34690 16322
rect 39678 16270 39730 16322
rect 2494 16158 2546 16210
rect 4622 16158 4674 16210
rect 7534 16158 7586 16210
rect 8542 16158 8594 16210
rect 16494 16158 16546 16210
rect 17054 16158 17106 16210
rect 17614 16158 17666 16210
rect 22430 16158 22482 16210
rect 22878 16158 22930 16210
rect 25566 16158 25618 16210
rect 38334 16158 38386 16210
rect 1822 16046 1874 16098
rect 5966 16046 6018 16098
rect 6414 16046 6466 16098
rect 7870 16046 7922 16098
rect 8094 16046 8146 16098
rect 9438 16046 9490 16098
rect 18958 16046 19010 16098
rect 25118 16046 25170 16098
rect 31614 16046 31666 16098
rect 34302 16046 34354 16098
rect 34526 16046 34578 16098
rect 37326 16046 37378 16098
rect 38894 16046 38946 16098
rect 7646 15934 7698 15986
rect 18286 15934 18338 15986
rect 22094 15934 22146 15986
rect 22318 15934 22370 15986
rect 23438 15934 23490 15986
rect 24334 15934 24386 15986
rect 24670 15934 24722 15986
rect 31950 15934 32002 15986
rect 33742 15934 33794 15986
rect 5070 15822 5122 15874
rect 6974 15822 7026 15874
rect 7534 15822 7586 15874
rect 9774 15822 9826 15874
rect 18062 15822 18114 15874
rect 19294 15822 19346 15874
rect 23326 15822 23378 15874
rect 33182 15822 33234 15874
rect 34638 15822 34690 15874
rect 36430 15822 36482 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 5630 15486 5682 15538
rect 6190 15486 6242 15538
rect 7758 15486 7810 15538
rect 9774 15486 9826 15538
rect 10782 15486 10834 15538
rect 16382 15486 16434 15538
rect 16830 15486 16882 15538
rect 17950 15486 18002 15538
rect 19742 15486 19794 15538
rect 29822 15486 29874 15538
rect 33406 15486 33458 15538
rect 37326 15486 37378 15538
rect 38894 15486 38946 15538
rect 39678 15486 39730 15538
rect 7646 15374 7698 15426
rect 8430 15374 8482 15426
rect 8990 15374 9042 15426
rect 11902 15374 11954 15426
rect 13694 15374 13746 15426
rect 14478 15374 14530 15426
rect 17726 15374 17778 15426
rect 18174 15374 18226 15426
rect 22542 15374 22594 15426
rect 25678 15374 25730 15426
rect 27246 15374 27298 15426
rect 29934 15374 29986 15426
rect 31614 15374 31666 15426
rect 33070 15374 33122 15426
rect 5518 15262 5570 15314
rect 6078 15262 6130 15314
rect 7198 15262 7250 15314
rect 7870 15262 7922 15314
rect 8766 15262 8818 15314
rect 9662 15262 9714 15314
rect 9886 15262 9938 15314
rect 10334 15262 10386 15314
rect 11566 15262 11618 15314
rect 13918 15262 13970 15314
rect 18510 15262 18562 15314
rect 19070 15262 19122 15314
rect 19406 15262 19458 15314
rect 19630 15262 19682 15314
rect 19854 15262 19906 15314
rect 19966 15262 20018 15314
rect 21870 15262 21922 15314
rect 30158 15262 30210 15314
rect 30494 15262 30546 15314
rect 30942 15262 30994 15314
rect 31166 15262 31218 15314
rect 31390 15262 31442 15314
rect 32174 15262 32226 15314
rect 8542 15150 8594 15202
rect 15374 15150 15426 15202
rect 18958 15150 19010 15202
rect 24670 15150 24722 15202
rect 25342 15150 25394 15202
rect 27470 15150 27522 15202
rect 38110 15150 38162 15202
rect 5630 15038 5682 15090
rect 6190 15038 6242 15090
rect 14366 15038 14418 15090
rect 18062 15038 18114 15090
rect 18734 15038 18786 15090
rect 31054 15038 31106 15090
rect 32174 15038 32226 15090
rect 32510 15038 32562 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16046 14702 16098 14754
rect 16718 14702 16770 14754
rect 18734 14702 18786 14754
rect 4958 14590 5010 14642
rect 5070 14590 5122 14642
rect 6190 14590 6242 14642
rect 7086 14590 7138 14642
rect 14590 14590 14642 14642
rect 17838 14590 17890 14642
rect 21422 14590 21474 14642
rect 23886 14590 23938 14642
rect 29150 14590 29202 14642
rect 30830 14590 30882 14642
rect 39566 14590 39618 14642
rect 5966 14478 6018 14530
rect 6974 14478 7026 14530
rect 12238 14478 12290 14530
rect 12350 14478 12402 14530
rect 12462 14478 12514 14530
rect 12574 14478 12626 14530
rect 12910 14478 12962 14530
rect 14030 14478 14082 14530
rect 14478 14478 14530 14530
rect 15710 14478 15762 14530
rect 18398 14478 18450 14530
rect 18958 14478 19010 14530
rect 19294 14478 19346 14530
rect 20078 14478 20130 14530
rect 20750 14478 20802 14530
rect 22206 14478 22258 14530
rect 22766 14478 22818 14530
rect 23438 14478 23490 14530
rect 23774 14478 23826 14530
rect 23998 14478 24050 14530
rect 25118 14478 25170 14530
rect 25902 14478 25954 14530
rect 29822 14478 29874 14530
rect 30046 14478 30098 14530
rect 31166 14478 31218 14530
rect 38894 14478 38946 14530
rect 4846 14366 4898 14418
rect 6638 14366 6690 14418
rect 13470 14366 13522 14418
rect 15038 14366 15090 14418
rect 15374 14366 15426 14418
rect 16158 14366 16210 14418
rect 16830 14366 16882 14418
rect 17390 14366 17442 14418
rect 17950 14366 18002 14418
rect 19742 14366 19794 14418
rect 24782 14366 24834 14418
rect 26574 14366 26626 14418
rect 36206 14366 36258 14418
rect 15598 14254 15650 14306
rect 16718 14254 16770 14306
rect 17614 14254 17666 14306
rect 17838 14254 17890 14306
rect 18622 14254 18674 14306
rect 19182 14254 19234 14306
rect 20414 14254 20466 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 5070 13918 5122 13970
rect 6078 13918 6130 13970
rect 8094 13918 8146 13970
rect 8206 13918 8258 13970
rect 8430 13918 8482 13970
rect 9662 13918 9714 13970
rect 13470 13918 13522 13970
rect 15486 13918 15538 13970
rect 18286 13918 18338 13970
rect 19406 13918 19458 13970
rect 20302 13918 20354 13970
rect 20750 13918 20802 13970
rect 25342 13918 25394 13970
rect 25454 13918 25506 13970
rect 28590 13918 28642 13970
rect 29822 13918 29874 13970
rect 30494 13918 30546 13970
rect 30718 13918 30770 13970
rect 2494 13806 2546 13858
rect 5742 13806 5794 13858
rect 5854 13806 5906 13858
rect 7534 13806 7586 13858
rect 7870 13806 7922 13858
rect 9998 13806 10050 13858
rect 11566 13806 11618 13858
rect 12238 13806 12290 13858
rect 16382 13806 16434 13858
rect 16830 13806 16882 13858
rect 17950 13806 18002 13858
rect 18174 13806 18226 13858
rect 19070 13806 19122 13858
rect 19182 13806 19234 13858
rect 25678 13806 25730 13858
rect 26910 13806 26962 13858
rect 30158 13806 30210 13858
rect 32174 13806 32226 13858
rect 35646 13806 35698 13858
rect 1822 13694 1874 13746
rect 8654 13694 8706 13746
rect 10334 13694 10386 13746
rect 11454 13694 11506 13746
rect 12014 13694 12066 13746
rect 12910 13694 12962 13746
rect 14030 13694 14082 13746
rect 15038 13694 15090 13746
rect 15598 13694 15650 13746
rect 15934 13694 15986 13746
rect 16606 13694 16658 13746
rect 17726 13694 17778 13746
rect 19854 13694 19906 13746
rect 25230 13694 25282 13746
rect 27470 13694 27522 13746
rect 28142 13694 28194 13746
rect 31166 13694 31218 13746
rect 31390 13694 31442 13746
rect 31614 13694 31666 13746
rect 32510 13694 32562 13746
rect 36430 13694 36482 13746
rect 4622 13582 4674 13634
rect 8318 13582 8370 13634
rect 13806 13582 13858 13634
rect 14702 13582 14754 13634
rect 15262 13582 15314 13634
rect 15486 13582 15538 13634
rect 16718 13582 16770 13634
rect 31838 13582 31890 13634
rect 33182 13582 33234 13634
rect 33518 13582 33570 13634
rect 36878 13582 36930 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 5742 13134 5794 13186
rect 7422 13134 7474 13186
rect 26686 13134 26738 13186
rect 27246 13134 27298 13186
rect 32286 13134 32338 13186
rect 32846 13134 32898 13186
rect 33070 13134 33122 13186
rect 7646 13022 7698 13074
rect 9662 13022 9714 13074
rect 33518 13022 33570 13074
rect 5518 12910 5570 12962
rect 8654 12910 8706 12962
rect 9214 12910 9266 12962
rect 9550 12910 9602 12962
rect 9998 12910 10050 12962
rect 10670 12910 10722 12962
rect 18734 12910 18786 12962
rect 19070 12910 19122 12962
rect 19518 12910 19570 12962
rect 21198 12910 21250 12962
rect 21534 12910 21586 12962
rect 21870 12910 21922 12962
rect 26350 12910 26402 12962
rect 30718 12910 30770 12962
rect 30830 12910 30882 12962
rect 31054 12910 31106 12962
rect 31278 12910 31330 12962
rect 31502 12910 31554 12962
rect 31838 12910 31890 12962
rect 32622 12910 32674 12962
rect 36430 12910 36482 12962
rect 38894 12910 38946 12962
rect 9886 12798 9938 12850
rect 10446 12798 10498 12850
rect 11790 12798 11842 12850
rect 13918 12798 13970 12850
rect 25566 12798 25618 12850
rect 26014 12798 26066 12850
rect 27134 12798 27186 12850
rect 30270 12798 30322 12850
rect 31726 12798 31778 12850
rect 35646 12798 35698 12850
rect 40014 12798 40066 12850
rect 5854 12686 5906 12738
rect 6078 12686 6130 12738
rect 7870 12686 7922 12738
rect 7982 12686 8034 12738
rect 8094 12686 8146 12738
rect 8766 12686 8818 12738
rect 8878 12686 8930 12738
rect 8990 12686 9042 12738
rect 11902 12686 11954 12738
rect 19294 12686 19346 12738
rect 19406 12686 19458 12738
rect 19630 12686 19682 12738
rect 21422 12686 21474 12738
rect 29934 12686 29986 12738
rect 32734 12686 32786 12738
rect 37102 12686 37154 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 6302 12350 6354 12402
rect 6638 12350 6690 12402
rect 8430 12350 8482 12402
rect 9550 12350 9602 12402
rect 9774 12350 9826 12402
rect 9998 12350 10050 12402
rect 11230 12350 11282 12402
rect 11566 12350 11618 12402
rect 13582 12350 13634 12402
rect 13694 12350 13746 12402
rect 13806 12350 13858 12402
rect 14926 12350 14978 12402
rect 18958 12350 19010 12402
rect 20526 12350 20578 12402
rect 25454 12350 25506 12402
rect 27918 12350 27970 12402
rect 31838 12350 31890 12402
rect 32286 12350 32338 12402
rect 33182 12350 33234 12402
rect 15934 12238 15986 12290
rect 16382 12238 16434 12290
rect 17614 12238 17666 12290
rect 20638 12238 20690 12290
rect 30942 12238 30994 12290
rect 31166 12238 31218 12290
rect 34078 12238 34130 12290
rect 40126 12238 40178 12290
rect 4846 12126 4898 12178
rect 5294 12126 5346 12178
rect 5742 12126 5794 12178
rect 7870 12126 7922 12178
rect 14254 12126 14306 12178
rect 14590 12126 14642 12178
rect 15710 12126 15762 12178
rect 17390 12126 17442 12178
rect 17838 12126 17890 12178
rect 17950 12126 18002 12178
rect 20078 12126 20130 12178
rect 20414 12126 20466 12178
rect 28030 12126 28082 12178
rect 28590 12126 28642 12178
rect 30830 12126 30882 12178
rect 31614 12126 31666 12178
rect 33630 12126 33682 12178
rect 33742 12126 33794 12178
rect 33966 12126 34018 12178
rect 4510 12014 4562 12066
rect 8094 12014 8146 12066
rect 9662 12014 9714 12066
rect 14030 12014 14082 12066
rect 16494 12014 16546 12066
rect 16606 12014 16658 12066
rect 17502 12014 17554 12066
rect 21086 12014 21138 12066
rect 5070 11902 5122 11954
rect 25230 11902 25282 11954
rect 25566 11902 25618 11954
rect 27918 11902 27970 11954
rect 28702 11902 28754 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 17614 11566 17666 11618
rect 19854 11566 19906 11618
rect 4846 11454 4898 11506
rect 9214 11454 9266 11506
rect 10558 11454 10610 11506
rect 13470 11454 13522 11506
rect 15150 11454 15202 11506
rect 18622 11454 18674 11506
rect 23214 11454 23266 11506
rect 25118 11454 25170 11506
rect 33854 11454 33906 11506
rect 2046 11342 2098 11394
rect 5630 11342 5682 11394
rect 6750 11342 6802 11394
rect 7198 11342 7250 11394
rect 7982 11342 8034 11394
rect 8430 11342 8482 11394
rect 8766 11342 8818 11394
rect 9438 11342 9490 11394
rect 9774 11342 9826 11394
rect 13582 11342 13634 11394
rect 14142 11342 14194 11394
rect 16830 11342 16882 11394
rect 17166 11342 17218 11394
rect 17614 11342 17666 11394
rect 17838 11342 17890 11394
rect 18174 11342 18226 11394
rect 20190 11342 20242 11394
rect 20414 11342 20466 11394
rect 21534 11342 21586 11394
rect 24446 11342 24498 11394
rect 25006 11342 25058 11394
rect 29150 11342 29202 11394
rect 32958 11342 33010 11394
rect 2718 11230 2770 11282
rect 5966 11230 6018 11282
rect 7646 11230 7698 11282
rect 8206 11230 8258 11282
rect 10110 11230 10162 11282
rect 16942 11230 16994 11282
rect 18958 11230 19010 11282
rect 21310 11230 21362 11282
rect 28142 11230 28194 11282
rect 28254 11230 28306 11282
rect 29486 11230 29538 11282
rect 33294 11230 33346 11282
rect 8766 11118 8818 11170
rect 9662 11118 9714 11170
rect 17390 11118 17442 11170
rect 19294 11118 19346 11170
rect 19966 11118 20018 11170
rect 27918 11118 27970 11170
rect 29262 11118 29314 11170
rect 31950 11118 32002 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 5854 10782 5906 10834
rect 6302 10782 6354 10834
rect 7534 10782 7586 10834
rect 8318 10782 8370 10834
rect 8766 10782 8818 10834
rect 11902 10782 11954 10834
rect 7646 10670 7698 10722
rect 8206 10670 8258 10722
rect 8542 10670 8594 10722
rect 12350 10782 12402 10834
rect 25454 10782 25506 10834
rect 27582 10782 27634 10834
rect 29934 10782 29986 10834
rect 10558 10670 10610 10722
rect 19630 10670 19682 10722
rect 24334 10670 24386 10722
rect 28926 10670 28978 10722
rect 2382 10558 2434 10610
rect 3054 10558 3106 10610
rect 5518 10558 5570 10610
rect 7310 10558 7362 10610
rect 8430 10558 8482 10610
rect 9662 10558 9714 10610
rect 9774 10558 9826 10610
rect 9998 10558 10050 10610
rect 10110 10558 10162 10610
rect 12126 10558 12178 10610
rect 12574 10558 12626 10610
rect 12910 10558 12962 10610
rect 22990 10558 23042 10610
rect 23662 10558 23714 10610
rect 24222 10558 24274 10610
rect 25342 10558 25394 10610
rect 25566 10558 25618 10610
rect 26014 10558 26066 10610
rect 27918 10558 27970 10610
rect 28590 10558 28642 10610
rect 29710 10558 29762 10610
rect 30046 10558 30098 10610
rect 30270 10558 30322 10610
rect 36430 10558 36482 10610
rect 36878 10558 36930 10610
rect 5182 10446 5234 10498
rect 8878 10446 8930 10498
rect 12238 10446 12290 10498
rect 13358 10446 13410 10498
rect 33518 10446 33570 10498
rect 35646 10446 35698 10498
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 8654 9998 8706 10050
rect 21422 9998 21474 10050
rect 29150 9998 29202 10050
rect 29486 9998 29538 10050
rect 12126 9886 12178 9938
rect 14030 9886 14082 9938
rect 16046 9886 16098 9938
rect 18174 9886 18226 9938
rect 18622 9886 18674 9938
rect 20526 9886 20578 9938
rect 20750 9886 20802 9938
rect 22318 9886 22370 9938
rect 23662 9886 23714 9938
rect 24782 9886 24834 9938
rect 25342 9886 25394 9938
rect 30942 9886 30994 9938
rect 31390 9886 31442 9938
rect 32846 9886 32898 9938
rect 34078 9886 34130 9938
rect 34862 9886 34914 9938
rect 8990 9774 9042 9826
rect 15374 9774 15426 9826
rect 21758 9774 21810 9826
rect 22206 9774 22258 9826
rect 23214 9774 23266 9826
rect 23438 9774 23490 9826
rect 23886 9774 23938 9826
rect 24222 9774 24274 9826
rect 26910 9774 26962 9826
rect 27806 9774 27858 9826
rect 32622 9774 32674 9826
rect 33854 9774 33906 9826
rect 34190 9774 34242 9826
rect 19070 9662 19122 9714
rect 19742 9662 19794 9714
rect 21310 9662 21362 9714
rect 24782 9662 24834 9714
rect 26350 9662 26402 9714
rect 29374 9662 29426 9714
rect 33294 9662 33346 9714
rect 34526 9662 34578 9714
rect 34750 9662 34802 9714
rect 8766 9550 8818 9602
rect 9438 9550 9490 9602
rect 12014 9550 12066 9602
rect 20078 9550 20130 9602
rect 21982 9550 22034 9602
rect 22318 9550 22370 9602
rect 22878 9550 22930 9602
rect 24446 9550 24498 9602
rect 24670 9550 24722 9602
rect 25230 9550 25282 9602
rect 27918 9550 27970 9602
rect 30382 9550 30434 9602
rect 31950 9550 32002 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 24558 9214 24610 9266
rect 25678 9214 25730 9266
rect 26014 9214 26066 9266
rect 26238 9214 26290 9266
rect 28142 9214 28194 9266
rect 28254 9214 28306 9266
rect 29150 9214 29202 9266
rect 11678 9102 11730 9154
rect 18734 9102 18786 9154
rect 18958 9102 19010 9154
rect 20638 9102 20690 9154
rect 23774 9102 23826 9154
rect 23886 9102 23938 9154
rect 25230 9102 25282 9154
rect 25454 9102 25506 9154
rect 27806 9102 27858 9154
rect 28590 9102 28642 9154
rect 31726 9102 31778 9154
rect 35198 9102 35250 9154
rect 10894 8990 10946 9042
rect 14926 8990 14978 9042
rect 19294 8990 19346 9042
rect 19406 8990 19458 9042
rect 19854 8990 19906 9042
rect 24334 8990 24386 9042
rect 24670 8990 24722 9042
rect 25902 8990 25954 9042
rect 26350 8990 26402 9042
rect 27134 8990 27186 9042
rect 27694 8990 27746 9042
rect 28366 8990 28418 9042
rect 32510 8990 32562 9042
rect 35870 8990 35922 9042
rect 36430 8990 36482 9042
rect 13806 8878 13858 8930
rect 14254 8878 14306 8930
rect 14702 8878 14754 8930
rect 19070 8878 19122 8930
rect 22766 8878 22818 8930
rect 29598 8878 29650 8930
rect 33070 8878 33122 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 14590 8430 14642 8482
rect 28366 8430 28418 8482
rect 32286 8430 32338 8482
rect 8878 8318 8930 8370
rect 11006 8318 11058 8370
rect 11454 8318 11506 8370
rect 14254 8318 14306 8370
rect 17054 8318 17106 8370
rect 19182 8318 19234 8370
rect 20078 8318 20130 8370
rect 20302 8318 20354 8370
rect 26126 8318 26178 8370
rect 27806 8318 27858 8370
rect 32398 8318 32450 8370
rect 8094 8206 8146 8258
rect 16382 8206 16434 8258
rect 19966 8206 20018 8258
rect 20526 8206 20578 8258
rect 21646 8206 21698 8258
rect 22094 8206 22146 8258
rect 27582 8206 27634 8258
rect 27918 8206 27970 8258
rect 28254 8206 28306 8258
rect 38894 8206 38946 8258
rect 14030 8094 14082 8146
rect 21422 8094 21474 8146
rect 21534 8094 21586 8146
rect 22766 8094 22818 8146
rect 40014 8094 40066 8146
rect 14366 7982 14418 8034
rect 15038 7982 15090 8034
rect 19742 7982 19794 8034
rect 22430 7982 22482 8034
rect 28366 7982 28418 8034
rect 32846 7982 32898 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 21086 7646 21138 7698
rect 40126 7646 40178 7698
rect 13918 7534 13970 7586
rect 39678 7534 39730 7586
rect 13134 7422 13186 7474
rect 16494 7422 16546 7474
rect 16046 7310 16098 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 25566 6862 25618 6914
rect 25230 6750 25282 6802
rect 21310 6638 21362 6690
rect 21534 6638 21586 6690
rect 21870 6638 21922 6690
rect 22318 6638 22370 6690
rect 26462 6638 26514 6690
rect 27470 6638 27522 6690
rect 22542 6526 22594 6578
rect 22990 6526 23042 6578
rect 24222 6526 24274 6578
rect 24334 6526 24386 6578
rect 24894 6526 24946 6578
rect 25454 6526 25506 6578
rect 26014 6526 26066 6578
rect 1710 6414 1762 6466
rect 21422 6414 21474 6466
rect 24558 6414 24610 6466
rect 25902 6414 25954 6466
rect 27134 6414 27186 6466
rect 40126 6414 40178 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 23214 6078 23266 6130
rect 1710 5966 1762 6018
rect 19518 5966 19570 6018
rect 23438 5966 23490 6018
rect 24670 5966 24722 6018
rect 26238 5966 26290 6018
rect 39790 5966 39842 6018
rect 18846 5854 18898 5906
rect 21982 5854 22034 5906
rect 22206 5854 22258 5906
rect 23102 5854 23154 5906
rect 24110 5854 24162 5906
rect 25566 5854 25618 5906
rect 28814 5854 28866 5906
rect 39566 5854 39618 5906
rect 40126 5854 40178 5906
rect 21646 5742 21698 5794
rect 24222 5742 24274 5794
rect 28366 5742 28418 5794
rect 22542 5630 22594 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 21310 5294 21362 5346
rect 26126 5294 26178 5346
rect 25790 5182 25842 5234
rect 21646 5070 21698 5122
rect 22878 5070 22930 5122
rect 26238 5070 26290 5122
rect 26462 5070 26514 5122
rect 38446 5070 38498 5122
rect 23662 4958 23714 5010
rect 38670 4958 38722 5010
rect 1710 4846 1762 4898
rect 21422 4846 21474 4898
rect 40126 4846 40178 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 24110 4510 24162 4562
rect 1710 4398 1762 4450
rect 20190 4398 20242 4450
rect 24334 4398 24386 4450
rect 39678 4398 39730 4450
rect 40126 4398 40178 4450
rect 19518 4286 19570 4338
rect 22318 4174 22370 4226
rect 23998 4174 24050 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 21198 3614 21250 3666
rect 20750 3502 20802 3554
rect 19630 3390 19682 3442
rect 19854 3390 19906 3442
rect 20190 3390 20242 3442
rect 1710 3278 1762 3330
rect 10334 3278 10386 3330
rect 11006 3278 11058 3330
rect 33182 3278 33234 3330
rect 39230 3278 39282 3330
rect 40126 3278 40178 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 8064 44685 8176 45485
rect 35616 44685 35728 45485
rect 8092 43708 8148 44685
rect 35644 43708 35700 44685
rect 8092 43652 8372 43708
rect 35644 43652 36036 43708
rect 8316 42194 8372 43652
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 8316 42142 8318 42194
rect 8370 42142 8372 42194
rect 8316 42130 8372 42142
rect 35980 42194 36036 43652
rect 35980 42142 35982 42194
rect 36034 42142 36036 42194
rect 35980 42130 36036 42142
rect 38780 43092 38836 43102
rect 38780 42194 38836 43036
rect 38780 42142 38782 42194
rect 38834 42142 38836 42194
rect 38780 42130 38836 42142
rect 40124 42420 40180 42430
rect 40124 42194 40180 42364
rect 40124 42142 40126 42194
rect 40178 42142 40180 42194
rect 40124 42130 40180 42142
rect 39228 42082 39284 42094
rect 39228 42030 39230 42082
rect 39282 42030 39284 42082
rect 39228 41748 39284 42030
rect 39228 41682 39284 41692
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 39676 41076 39732 41086
rect 39676 40982 39732 41020
rect 1708 40962 1764 40974
rect 1708 40910 1710 40962
rect 1762 40910 1764 40962
rect 1708 40404 1764 40910
rect 29372 40962 29428 40974
rect 30380 40964 30436 40974
rect 29372 40910 29374 40962
rect 29426 40910 29428 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 1708 40338 1764 40348
rect 25900 40404 25956 40414
rect 25900 40310 25956 40348
rect 26796 40404 26852 40414
rect 26572 40292 26628 40302
rect 26572 40198 26628 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4284 39732 4340 39742
rect 26348 39732 26404 39742
rect 1708 37378 1764 37390
rect 1708 37326 1710 37378
rect 1762 37326 1764 37378
rect 1708 37044 1764 37326
rect 1708 36978 1764 36988
rect 1708 36372 1764 36382
rect 1708 36278 1764 36316
rect 3948 26964 4004 26974
rect 2044 26402 2100 26414
rect 2044 26350 2046 26402
rect 2098 26350 2100 26402
rect 1820 26290 1876 26302
rect 1820 26238 1822 26290
rect 1874 26238 1876 26290
rect 1708 25618 1764 25630
rect 1708 25566 1710 25618
rect 1762 25566 1764 25618
rect 1708 25172 1764 25566
rect 1708 25106 1764 25116
rect 1708 24948 1764 24958
rect 1820 24948 1876 26238
rect 2044 25396 2100 26350
rect 3948 26402 4004 26908
rect 3948 26350 3950 26402
rect 4002 26350 4004 26402
rect 2044 25330 2100 25340
rect 2492 26178 2548 26190
rect 2492 26126 2494 26178
rect 2546 26126 2548 26178
rect 1764 24892 1876 24948
rect 2492 24948 2548 26126
rect 3836 26066 3892 26078
rect 3836 26014 3838 26066
rect 3890 26014 3892 26066
rect 3836 25618 3892 26014
rect 3836 25566 3838 25618
rect 3890 25566 3892 25618
rect 3836 25554 3892 25566
rect 2940 25172 2996 25182
rect 1708 24882 1764 24892
rect 2492 24882 2548 24892
rect 2828 25116 2940 25172
rect 1708 24610 1764 24622
rect 1708 24558 1710 24610
rect 1762 24558 1764 24610
rect 1708 21812 1764 24558
rect 1932 24276 1988 24286
rect 1932 24050 1988 24220
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23986 1988 23998
rect 1708 21746 1764 21756
rect 2828 21700 2884 25116
rect 2940 25106 2996 25116
rect 3836 24610 3892 24622
rect 3836 24558 3838 24610
rect 3890 24558 3892 24610
rect 2940 24164 2996 24174
rect 2940 23938 2996 24108
rect 3836 24162 3892 24558
rect 3836 24110 3838 24162
rect 3890 24110 3892 24162
rect 3836 24098 3892 24110
rect 2940 23886 2942 23938
rect 2994 23886 2996 23938
rect 2940 23874 2996 23886
rect 3836 23940 3892 23950
rect 3948 23940 4004 26350
rect 4172 26066 4228 26078
rect 4172 26014 4174 26066
rect 4226 26014 4228 26066
rect 4172 25060 4228 26014
rect 4172 24994 4228 25004
rect 4172 24612 4228 24622
rect 4172 24162 4228 24556
rect 4172 24110 4174 24162
rect 4226 24110 4228 24162
rect 4172 24098 4228 24110
rect 3836 23938 4004 23940
rect 3836 23886 3838 23938
rect 3890 23886 4004 23938
rect 3836 23884 4004 23886
rect 3276 23380 3332 23390
rect 3052 21812 3108 21822
rect 3052 21718 3108 21756
rect 2940 21700 2996 21710
rect 2716 21698 2996 21700
rect 2716 21646 2942 21698
rect 2994 21646 2996 21698
rect 2716 21644 2996 21646
rect 1708 20690 1764 20702
rect 1708 20638 1710 20690
rect 1762 20638 1764 20690
rect 1708 20244 1764 20638
rect 1708 20178 1764 20188
rect 2044 20578 2100 20590
rect 2044 20526 2046 20578
rect 2098 20526 2100 20578
rect 2044 20020 2100 20526
rect 2380 20580 2436 20590
rect 2380 20242 2436 20524
rect 2380 20190 2382 20242
rect 2434 20190 2436 20242
rect 2380 20178 2436 20190
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 2492 20244 2548 20526
rect 2492 20178 2548 20188
rect 2156 20020 2212 20030
rect 1932 20018 2212 20020
rect 1932 19966 2158 20018
rect 2210 19966 2212 20018
rect 1932 19964 2212 19966
rect 1708 19572 1764 19582
rect 1708 19234 1764 19516
rect 1708 19182 1710 19234
rect 1762 19182 1764 19234
rect 1708 19170 1764 19182
rect 1932 18452 1988 19964
rect 2156 19954 2212 19964
rect 2716 20020 2772 21644
rect 2940 21634 2996 21644
rect 3052 21364 3108 21374
rect 2716 19926 2772 19964
rect 2828 21362 3108 21364
rect 2828 21310 3054 21362
rect 3106 21310 3108 21362
rect 2828 21308 3108 21310
rect 2492 19572 2548 19582
rect 2492 19346 2548 19516
rect 2492 19294 2494 19346
rect 2546 19294 2548 19346
rect 2492 19282 2548 19294
rect 2828 19348 2884 21308
rect 3052 21298 3108 21308
rect 3164 20690 3220 20702
rect 3164 20638 3166 20690
rect 3218 20638 3220 20690
rect 2828 19282 2884 19292
rect 2940 20578 2996 20590
rect 2940 20526 2942 20578
rect 2994 20526 2996 20578
rect 2940 19348 2996 20526
rect 3052 20578 3108 20590
rect 3052 20526 3054 20578
rect 3106 20526 3108 20578
rect 3052 19908 3108 20526
rect 3052 19842 3108 19852
rect 3164 20244 3220 20638
rect 3276 20468 3332 23324
rect 3836 23380 3892 23884
rect 3836 23314 3892 23324
rect 4284 23044 4340 39676
rect 26124 39730 26404 39732
rect 26124 39678 26350 39730
rect 26402 39678 26404 39730
rect 26124 39676 26404 39678
rect 23548 39618 23604 39630
rect 23548 39566 23550 39618
rect 23602 39566 23604 39618
rect 23548 39396 23604 39566
rect 24220 39508 24276 39518
rect 24220 39414 24276 39452
rect 25340 39508 25396 39518
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 11340 38836 11396 38846
rect 23212 38836 23268 38846
rect 11340 38834 11508 38836
rect 11340 38782 11342 38834
rect 11394 38782 11508 38834
rect 11340 38780 11508 38782
rect 11340 38770 11396 38780
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 8428 37828 8484 37838
rect 8204 37044 8260 37054
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 8204 36594 8260 36988
rect 8204 36542 8206 36594
rect 8258 36542 8260 36594
rect 8204 36530 8260 36542
rect 7532 36482 7588 36494
rect 7532 36430 7534 36482
rect 7586 36430 7588 36482
rect 6972 35588 7028 35598
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 5628 33460 5684 33470
rect 5628 33366 5684 33404
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5964 30324 6020 30334
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 5964 28866 6020 30268
rect 5964 28814 5966 28866
rect 6018 28814 6020 28866
rect 5964 28802 6020 28814
rect 5628 28756 5684 28766
rect 5404 28754 5684 28756
rect 5404 28702 5630 28754
rect 5682 28702 5684 28754
rect 5404 28700 5684 28702
rect 4732 28644 4788 28654
rect 4732 27860 4788 28588
rect 5404 27970 5460 28700
rect 5628 28690 5684 28700
rect 6300 28644 6356 28654
rect 6300 28550 6356 28588
rect 5740 28420 5796 28430
rect 5404 27918 5406 27970
rect 5458 27918 5460 27970
rect 5404 27906 5460 27918
rect 5628 28418 5796 28420
rect 5628 28366 5742 28418
rect 5794 28366 5796 28418
rect 5628 28364 5796 28366
rect 4732 27858 4900 27860
rect 4732 27806 4734 27858
rect 4786 27806 4900 27858
rect 4732 27804 4900 27806
rect 4732 27794 4788 27804
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4620 25508 4676 25518
rect 4844 25508 4900 27804
rect 5628 26964 5684 28364
rect 5740 28354 5796 28364
rect 6972 27300 7028 35532
rect 7532 33236 7588 36430
rect 8428 35924 8484 37772
rect 9660 37828 9716 37838
rect 9660 37490 9716 37772
rect 9660 37438 9662 37490
rect 9714 37438 9716 37490
rect 9660 37426 9716 37438
rect 9548 37044 9604 37054
rect 9548 36950 9604 36988
rect 9884 37042 9940 37054
rect 9884 36990 9886 37042
rect 9938 36990 9940 37042
rect 9884 36596 9940 36990
rect 9884 36530 9940 36540
rect 10332 36596 10388 36606
rect 10332 36594 10836 36596
rect 10332 36542 10334 36594
rect 10386 36542 10836 36594
rect 10332 36540 10836 36542
rect 10332 36530 10388 36540
rect 7868 35922 8484 35924
rect 7868 35870 8430 35922
rect 8482 35870 8484 35922
rect 7868 35868 8484 35870
rect 7868 34354 7924 35868
rect 8428 35858 8484 35868
rect 9772 36260 9828 36270
rect 9772 35810 9828 36204
rect 9996 35812 10052 35822
rect 9772 35758 9774 35810
rect 9826 35758 9828 35810
rect 9772 35746 9828 35758
rect 9884 35810 10052 35812
rect 9884 35758 9998 35810
rect 10050 35758 10052 35810
rect 9884 35756 10052 35758
rect 8204 35698 8260 35710
rect 8204 35646 8206 35698
rect 8258 35646 8260 35698
rect 8204 35588 8260 35646
rect 8204 35522 8260 35532
rect 8876 35588 8932 35598
rect 8876 35494 8932 35532
rect 7868 34302 7870 34354
rect 7922 34302 7924 34354
rect 7868 34290 7924 34302
rect 9772 34356 9828 34366
rect 9884 34356 9940 35756
rect 9996 35746 10052 35756
rect 10444 35812 10500 35822
rect 10220 34914 10276 34926
rect 10220 34862 10222 34914
rect 10274 34862 10276 34914
rect 10220 34692 10276 34862
rect 10444 34802 10500 35756
rect 10444 34750 10446 34802
rect 10498 34750 10500 34802
rect 10444 34738 10500 34750
rect 10780 35364 10836 36540
rect 10780 34914 10836 35308
rect 10780 34862 10782 34914
rect 10834 34862 10836 34914
rect 10220 34626 10276 34636
rect 10780 34468 10836 34862
rect 11228 35700 11284 35710
rect 11228 35026 11284 35644
rect 11228 34974 11230 35026
rect 11282 34974 11284 35026
rect 10780 34412 11172 34468
rect 9772 34354 9940 34356
rect 9772 34302 9774 34354
rect 9826 34302 9940 34354
rect 9772 34300 9940 34302
rect 10332 34300 10724 34356
rect 9772 34290 9828 34300
rect 8988 34242 9044 34254
rect 8988 34190 8990 34242
rect 9042 34190 9044 34242
rect 8764 34130 8820 34142
rect 8764 34078 8766 34130
rect 8818 34078 8820 34130
rect 7756 33906 7812 33918
rect 7756 33854 7758 33906
rect 7810 33854 7812 33906
rect 7756 33458 7812 33854
rect 7756 33406 7758 33458
rect 7810 33406 7812 33458
rect 7756 33394 7812 33406
rect 8092 33906 8148 33918
rect 8092 33854 8094 33906
rect 8146 33854 8148 33906
rect 7532 33170 7588 33180
rect 7644 32674 7700 32686
rect 7644 32622 7646 32674
rect 7698 32622 7700 32674
rect 7644 32564 7700 32622
rect 7644 30100 7700 32508
rect 7980 32562 8036 32574
rect 7980 32510 7982 32562
rect 8034 32510 8036 32562
rect 7980 31556 8036 32510
rect 8092 32452 8148 33854
rect 8764 33460 8820 34078
rect 8764 33394 8820 33404
rect 8540 33346 8596 33358
rect 8540 33294 8542 33346
rect 8594 33294 8596 33346
rect 8540 33236 8596 33294
rect 8876 33236 8932 33246
rect 8540 33170 8596 33180
rect 8652 33234 8932 33236
rect 8652 33182 8878 33234
rect 8930 33182 8932 33234
rect 8652 33180 8932 33182
rect 8540 32788 8596 32798
rect 8652 32788 8708 33180
rect 8876 33170 8932 33180
rect 8540 32786 8708 32788
rect 8540 32734 8542 32786
rect 8594 32734 8708 32786
rect 8540 32732 8708 32734
rect 8764 33012 8820 33022
rect 8988 33012 9044 34190
rect 9660 34132 9716 34142
rect 9660 34038 9716 34076
rect 9884 34130 9940 34142
rect 9884 34078 9886 34130
rect 9938 34078 9940 34130
rect 9212 34020 9268 34030
rect 9212 33460 9268 33964
rect 9884 33908 9940 34078
rect 10332 34130 10388 34300
rect 10332 34078 10334 34130
rect 10386 34078 10388 34130
rect 10332 34066 10388 34078
rect 10556 34130 10612 34142
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 10556 33908 10612 34078
rect 9548 33852 10612 33908
rect 9212 33458 9492 33460
rect 9212 33406 9214 33458
rect 9266 33406 9492 33458
rect 9212 33404 9492 33406
rect 9212 33394 9268 33404
rect 8820 32956 9044 33012
rect 8764 32786 8820 32956
rect 8764 32734 8766 32786
rect 8818 32734 8820 32786
rect 8540 32722 8596 32732
rect 8764 32722 8820 32734
rect 8316 32674 8372 32686
rect 8316 32622 8318 32674
rect 8370 32622 8372 32674
rect 8204 32564 8260 32574
rect 8316 32564 8372 32622
rect 8260 32508 8372 32564
rect 8988 32562 9044 32574
rect 8988 32510 8990 32562
rect 9042 32510 9044 32562
rect 8204 32498 8260 32508
rect 8092 32386 8148 32396
rect 8652 32452 8708 32462
rect 8652 32358 8708 32396
rect 8316 31556 8372 31566
rect 7980 31554 8372 31556
rect 7980 31502 8318 31554
rect 8370 31502 8372 31554
rect 7980 31500 8372 31502
rect 8316 31220 8372 31500
rect 8316 31154 8372 31164
rect 8988 31556 9044 32510
rect 9212 31556 9268 31566
rect 8988 31500 9212 31556
rect 8988 30436 9044 31500
rect 9212 31462 9268 31500
rect 8540 30380 9044 30436
rect 8204 30324 8260 30334
rect 8204 30230 8260 30268
rect 8540 30210 8596 30380
rect 8988 30322 9044 30380
rect 8988 30270 8990 30322
rect 9042 30270 9044 30322
rect 8988 30258 9044 30270
rect 8540 30158 8542 30210
rect 8594 30158 8596 30210
rect 8540 30146 8596 30158
rect 8876 30212 8932 30222
rect 7868 30100 7924 30110
rect 7644 30098 7924 30100
rect 7644 30046 7870 30098
rect 7922 30046 7924 30098
rect 7644 30044 7924 30046
rect 7532 29988 7588 29998
rect 7084 29316 7140 29326
rect 7084 28754 7140 29260
rect 7084 28702 7086 28754
rect 7138 28702 7140 28754
rect 7084 28690 7140 28702
rect 7532 27746 7588 29932
rect 7532 27694 7534 27746
rect 7586 27694 7588 27746
rect 7532 27682 7588 27694
rect 6972 27188 7028 27244
rect 6524 27186 7028 27188
rect 6524 27134 6974 27186
rect 7026 27134 7028 27186
rect 6524 27132 7028 27134
rect 6524 27074 6580 27132
rect 6972 27122 7028 27132
rect 6524 27022 6526 27074
rect 6578 27022 6580 27074
rect 6524 27010 6580 27022
rect 5628 26898 5684 26908
rect 6188 26964 6244 27002
rect 7868 26908 7924 30044
rect 8092 29986 8148 29998
rect 8092 29934 8094 29986
rect 8146 29934 8148 29986
rect 7980 29540 8036 29550
rect 8092 29540 8148 29934
rect 8316 29988 8372 29998
rect 8316 29894 8372 29932
rect 7980 29538 8148 29540
rect 7980 29486 7982 29538
rect 8034 29486 8148 29538
rect 7980 29484 8148 29486
rect 7980 29474 8036 29484
rect 8652 29428 8708 29438
rect 8652 29334 8708 29372
rect 8876 29426 8932 30156
rect 9436 29986 9492 33404
rect 9548 33346 9604 33852
rect 9548 33294 9550 33346
rect 9602 33294 9604 33346
rect 9548 33282 9604 33294
rect 9660 33460 9716 33470
rect 9660 32562 9716 33404
rect 10556 32674 10612 33852
rect 10668 33908 10724 34300
rect 10892 34244 10948 34254
rect 10668 33842 10724 33852
rect 10780 34188 10892 34244
rect 10668 33684 10724 33694
rect 10668 33234 10724 33628
rect 10668 33182 10670 33234
rect 10722 33182 10724 33234
rect 10668 33170 10724 33182
rect 10556 32622 10558 32674
rect 10610 32622 10612 32674
rect 10556 32610 10612 32622
rect 9660 32510 9662 32562
rect 9714 32510 9716 32562
rect 9660 32498 9716 32510
rect 10108 32562 10164 32574
rect 10108 32510 10110 32562
rect 10162 32510 10164 32562
rect 10108 32004 10164 32510
rect 10108 30994 10164 31948
rect 10108 30942 10110 30994
rect 10162 30942 10164 30994
rect 10108 30930 10164 30942
rect 9548 30770 9604 30782
rect 9548 30718 9550 30770
rect 9602 30718 9604 30770
rect 9548 30210 9604 30718
rect 9884 30772 9940 30782
rect 9884 30770 10052 30772
rect 9884 30718 9886 30770
rect 9938 30718 10052 30770
rect 9884 30716 10052 30718
rect 9884 30706 9940 30716
rect 9996 30324 10052 30716
rect 10780 30324 10836 34188
rect 10892 34178 10948 34188
rect 11004 34132 11060 34142
rect 10892 34020 10948 34030
rect 10892 33926 10948 33964
rect 11004 33458 11060 34076
rect 11004 33406 11006 33458
rect 11058 33406 11060 33458
rect 11004 33394 11060 33406
rect 11116 33346 11172 34412
rect 11116 33294 11118 33346
rect 11170 33294 11172 33346
rect 11116 33282 11172 33294
rect 10892 33122 10948 33134
rect 10892 33070 10894 33122
rect 10946 33070 10948 33122
rect 10892 33012 10948 33070
rect 11228 33012 11284 34974
rect 11340 33908 11396 33918
rect 11340 33346 11396 33852
rect 11340 33294 11342 33346
rect 11394 33294 11396 33346
rect 11340 33282 11396 33294
rect 11452 33236 11508 38780
rect 12012 38724 12068 38734
rect 14140 38724 14196 38734
rect 12012 38722 12404 38724
rect 12012 38670 12014 38722
rect 12066 38670 12404 38722
rect 12012 38668 12404 38670
rect 12012 38658 12068 38668
rect 12348 38274 12404 38668
rect 14140 38722 14308 38724
rect 14140 38670 14142 38722
rect 14194 38670 14308 38722
rect 14140 38668 14308 38670
rect 14140 38658 14196 38668
rect 12348 38222 12350 38274
rect 12402 38222 12404 38274
rect 12348 38210 12404 38222
rect 14252 38162 14308 38668
rect 14252 38110 14254 38162
rect 14306 38110 14308 38162
rect 14140 38050 14196 38062
rect 14140 37998 14142 38050
rect 14194 37998 14196 38050
rect 12684 37938 12740 37950
rect 12684 37886 12686 37938
rect 12738 37886 12740 37938
rect 12460 37828 12516 37838
rect 12460 37734 12516 37772
rect 12124 36596 12180 36606
rect 12124 36502 12180 36540
rect 12684 36596 12740 37886
rect 13468 37938 13524 37950
rect 13468 37886 13470 37938
rect 13522 37886 13524 37938
rect 13356 37828 13412 37838
rect 12684 36530 12740 36540
rect 13244 37380 13300 37390
rect 12012 36484 12068 36494
rect 12012 36390 12068 36428
rect 12684 36372 12740 36382
rect 12684 36278 12740 36316
rect 12236 36258 12292 36270
rect 12236 36206 12238 36258
rect 12290 36206 12292 36258
rect 11676 35812 11732 35822
rect 11676 35718 11732 35756
rect 12236 35700 12292 36206
rect 12460 36260 12516 36270
rect 12460 36166 12516 36204
rect 12236 35634 12292 35644
rect 11676 35364 11732 35374
rect 11676 35138 11732 35308
rect 11676 35086 11678 35138
rect 11730 35086 11732 35138
rect 11676 35074 11732 35086
rect 12012 34916 12068 34926
rect 13244 34916 13300 37324
rect 13356 36820 13412 37772
rect 13468 37492 13524 37886
rect 13692 37492 13748 37502
rect 13468 37436 13692 37492
rect 13468 37266 13524 37278
rect 13468 37214 13470 37266
rect 13522 37214 13524 37266
rect 13468 37044 13524 37214
rect 13580 37154 13636 37436
rect 13692 37426 13748 37436
rect 14140 37380 14196 37998
rect 14140 37314 14196 37324
rect 14252 37828 14308 38110
rect 16268 38162 16324 38174
rect 16268 38110 16270 38162
rect 16322 38110 16324 38162
rect 15484 37940 15540 37950
rect 15260 37938 15540 37940
rect 15260 37886 15486 37938
rect 15538 37886 15540 37938
rect 15260 37884 15540 37886
rect 14812 37828 14868 37838
rect 14252 37826 14868 37828
rect 14252 37774 14814 37826
rect 14866 37774 14868 37826
rect 14252 37772 14868 37774
rect 14028 37156 14084 37166
rect 13580 37102 13582 37154
rect 13634 37102 13636 37154
rect 13580 37090 13636 37102
rect 13692 37154 14084 37156
rect 13692 37102 14030 37154
rect 14082 37102 14084 37154
rect 13692 37100 14084 37102
rect 13468 36978 13524 36988
rect 13356 36764 13524 36820
rect 13468 36148 13524 36764
rect 13580 36482 13636 36494
rect 13580 36430 13582 36482
rect 13634 36430 13636 36482
rect 13580 36372 13636 36430
rect 13692 36482 13748 37100
rect 14028 37090 14084 37100
rect 13804 36596 13860 36606
rect 13804 36502 13860 36540
rect 13692 36430 13694 36482
rect 13746 36430 13748 36482
rect 13692 36418 13748 36430
rect 14028 36484 14084 36494
rect 14028 36390 14084 36428
rect 13580 36306 13636 36316
rect 13916 36260 13972 36270
rect 13916 36166 13972 36204
rect 13468 36092 13636 36148
rect 13468 35586 13524 35598
rect 13468 35534 13470 35586
rect 13522 35534 13524 35586
rect 13468 35364 13524 35534
rect 13580 35476 13636 36092
rect 13692 35700 13748 35710
rect 14252 35700 14308 37772
rect 14812 37762 14868 37772
rect 15148 37826 15204 37838
rect 15148 37774 15150 37826
rect 15202 37774 15204 37826
rect 15148 37604 15204 37774
rect 15036 37548 15204 37604
rect 14812 37156 14868 37166
rect 14868 37100 14980 37156
rect 14812 37062 14868 37100
rect 14812 36932 14868 36942
rect 13692 35698 14308 35700
rect 13692 35646 13694 35698
rect 13746 35646 14308 35698
rect 13692 35644 14308 35646
rect 14588 36258 14644 36270
rect 14588 36206 14590 36258
rect 14642 36206 14644 36258
rect 13692 35634 13748 35644
rect 14028 35476 14084 35486
rect 13580 35420 13748 35476
rect 13468 35298 13524 35308
rect 12012 34914 13300 34916
rect 12012 34862 12014 34914
rect 12066 34862 13300 34914
rect 12012 34860 13300 34862
rect 12012 34850 12068 34860
rect 11452 33170 11508 33180
rect 11564 34692 11620 34702
rect 11564 33684 11620 34636
rect 11788 34690 11844 34702
rect 11788 34638 11790 34690
rect 11842 34638 11844 34690
rect 11788 34130 11844 34638
rect 12012 34580 12068 34590
rect 12012 34242 12068 34524
rect 12012 34190 12014 34242
rect 12066 34190 12068 34242
rect 12012 34178 12068 34190
rect 11788 34078 11790 34130
rect 11842 34078 11844 34130
rect 11788 34066 11844 34078
rect 12124 34132 12180 34142
rect 12124 34038 12180 34076
rect 11564 33234 11620 33628
rect 11564 33182 11566 33234
rect 11618 33182 11620 33234
rect 11564 33170 11620 33182
rect 11676 33234 11732 33246
rect 11676 33182 11678 33234
rect 11730 33182 11732 33234
rect 11676 33012 11732 33182
rect 11228 32956 11620 33012
rect 10892 32946 10948 32956
rect 11452 31668 11508 31678
rect 11452 30996 11508 31612
rect 11004 30994 11508 30996
rect 11004 30942 11454 30994
rect 11506 30942 11508 30994
rect 11004 30940 11508 30942
rect 10892 30324 10948 30334
rect 9996 30268 10164 30324
rect 9884 30212 9940 30222
rect 9548 30158 9550 30210
rect 9602 30158 9604 30210
rect 9548 30146 9604 30158
rect 9660 30156 9884 30212
rect 9436 29934 9438 29986
rect 9490 29934 9492 29986
rect 9436 29922 9492 29934
rect 9660 29652 9716 30156
rect 9884 30118 9940 30156
rect 9548 29596 9716 29652
rect 9996 30098 10052 30110
rect 9996 30046 9998 30098
rect 10050 30046 10052 30098
rect 8876 29374 8878 29426
rect 8930 29374 8932 29426
rect 8876 29362 8932 29374
rect 9436 29428 9492 29438
rect 9212 28756 9268 28766
rect 9212 28662 9268 28700
rect 9436 27636 9492 29372
rect 9548 28754 9604 29596
rect 9996 29540 10052 30046
rect 9884 29484 10052 29540
rect 10108 29988 10164 30268
rect 9660 29426 9716 29438
rect 9660 29374 9662 29426
rect 9714 29374 9716 29426
rect 9660 28868 9716 29374
rect 9772 29428 9828 29438
rect 9772 29334 9828 29372
rect 9660 28812 9828 28868
rect 9548 28702 9550 28754
rect 9602 28702 9604 28754
rect 9548 28690 9604 28702
rect 9660 28084 9716 28094
rect 9772 28084 9828 28812
rect 9884 28756 9940 29484
rect 9996 29316 10052 29326
rect 9996 29222 10052 29260
rect 10108 28980 10164 29932
rect 10220 30322 10948 30324
rect 10220 30270 10894 30322
rect 10946 30270 10948 30322
rect 10220 30268 10948 30270
rect 10220 29426 10276 30268
rect 10220 29374 10222 29426
rect 10274 29374 10276 29426
rect 10220 29362 10276 29374
rect 10108 28914 10164 28924
rect 10332 29204 10388 29214
rect 9884 28690 9940 28700
rect 10220 28644 10276 28654
rect 10332 28644 10388 29148
rect 10444 28980 10500 28990
rect 10444 28754 10500 28924
rect 10444 28702 10446 28754
rect 10498 28702 10500 28754
rect 10444 28690 10500 28702
rect 10220 28642 10388 28644
rect 10220 28590 10222 28642
rect 10274 28590 10388 28642
rect 10220 28588 10388 28590
rect 10220 28578 10276 28588
rect 9660 28082 9828 28084
rect 9660 28030 9662 28082
rect 9714 28030 9828 28082
rect 9660 28028 9828 28030
rect 9660 28018 9716 28028
rect 9548 27860 9604 27870
rect 9548 27766 9604 27804
rect 9772 27858 9828 27870
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 9772 27636 9828 27806
rect 10220 27860 10276 27870
rect 10220 27858 10388 27860
rect 10220 27806 10222 27858
rect 10274 27806 10388 27858
rect 10220 27804 10388 27806
rect 10220 27794 10276 27804
rect 9436 27580 9828 27636
rect 6188 26898 6244 26908
rect 4620 25506 4900 25508
rect 4620 25454 4622 25506
rect 4674 25454 4900 25506
rect 4620 25452 4900 25454
rect 7308 26852 7924 26908
rect 9436 27412 9492 27422
rect 4620 24724 4676 25452
rect 4620 24630 4676 24668
rect 5068 25172 5124 25182
rect 5068 24722 5124 25116
rect 6412 25060 6468 25070
rect 6468 25004 6580 25060
rect 6412 24994 6468 25004
rect 6524 24946 6580 25004
rect 6524 24894 6526 24946
rect 6578 24894 6580 24946
rect 6524 24882 6580 24894
rect 5292 24836 5348 24846
rect 5292 24742 5348 24780
rect 6412 24836 6468 24846
rect 5068 24670 5070 24722
rect 5122 24670 5124 24722
rect 5068 24658 5124 24670
rect 6300 24722 6356 24734
rect 6300 24670 6302 24722
rect 6354 24670 6356 24722
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 6300 23940 6356 24670
rect 6412 24722 6468 24780
rect 6860 24836 6916 24846
rect 7308 24836 7364 26852
rect 6860 24834 7364 24836
rect 6860 24782 6862 24834
rect 6914 24782 7364 24834
rect 6860 24780 7364 24782
rect 6860 24770 6916 24780
rect 6412 24670 6414 24722
rect 6466 24670 6468 24722
rect 6412 24052 6468 24670
rect 6636 24722 6692 24734
rect 6636 24670 6638 24722
rect 6690 24670 6692 24722
rect 6636 24052 6692 24670
rect 7308 24722 7364 24780
rect 8652 25284 8708 25294
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 24658 7364 24670
rect 7420 24722 7476 24734
rect 7420 24670 7422 24722
rect 7474 24670 7476 24722
rect 6412 23996 6580 24052
rect 6636 23996 6804 24052
rect 6524 23940 6580 23996
rect 6524 23884 6692 23940
rect 6300 23874 6356 23884
rect 6412 23826 6468 23838
rect 6412 23774 6414 23826
rect 6466 23774 6468 23826
rect 4732 23716 4788 23726
rect 4732 23378 4788 23660
rect 5292 23492 5348 23502
rect 4732 23326 4734 23378
rect 4786 23326 4788 23378
rect 4732 23314 4788 23326
rect 5180 23380 5236 23390
rect 4508 23266 4564 23278
rect 4508 23214 4510 23266
rect 4562 23214 4564 23266
rect 4396 23156 4452 23166
rect 4396 23062 4452 23100
rect 4284 22978 4340 22988
rect 4508 22932 4564 23214
rect 5068 23268 5124 23278
rect 5068 23174 5124 23212
rect 4508 22866 4564 22876
rect 4956 23154 5012 23166
rect 4956 23102 4958 23154
rect 5010 23102 5012 23154
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4956 22596 5012 23102
rect 4956 22530 5012 22540
rect 5068 22484 5124 22494
rect 5068 22390 5124 22428
rect 4732 22370 4788 22382
rect 4732 22318 4734 22370
rect 4786 22318 4788 22370
rect 4732 22260 4788 22318
rect 4844 22260 4900 22270
rect 4732 22204 4844 22260
rect 4844 22194 4900 22204
rect 4956 22260 5012 22270
rect 5180 22260 5236 23324
rect 5292 23378 5348 23436
rect 5292 23326 5294 23378
rect 5346 23326 5348 23378
rect 5292 23314 5348 23326
rect 5964 23266 6020 23278
rect 5964 23214 5966 23266
rect 6018 23214 6020 23266
rect 5516 23156 5572 23166
rect 4956 22258 5236 22260
rect 4956 22206 4958 22258
rect 5010 22206 5236 22258
rect 4956 22204 5236 22206
rect 5292 23154 5572 23156
rect 5292 23102 5518 23154
rect 5570 23102 5572 23154
rect 5292 23100 5572 23102
rect 4956 22194 5012 22204
rect 3500 21812 3556 21822
rect 3500 21718 3556 21756
rect 4844 21812 4900 21822
rect 5068 21812 5124 22204
rect 4844 21810 5124 21812
rect 4844 21758 4846 21810
rect 4898 21758 5124 21810
rect 4844 21756 5124 21758
rect 4844 21746 4900 21756
rect 3836 21698 3892 21710
rect 3836 21646 3838 21698
rect 3890 21646 3892 21698
rect 3836 21588 3892 21646
rect 5068 21700 5124 21756
rect 5068 21634 5124 21644
rect 3836 21522 3892 21532
rect 4620 21588 4676 21598
rect 5180 21588 5236 21598
rect 5292 21588 5348 23100
rect 5516 23090 5572 23100
rect 5628 23156 5684 23166
rect 5628 23062 5684 23100
rect 5740 23154 5796 23166
rect 5740 23102 5742 23154
rect 5794 23102 5796 23154
rect 5628 22820 5684 22830
rect 5516 22708 5572 22718
rect 5404 22148 5460 22158
rect 5404 21810 5460 22092
rect 5404 21758 5406 21810
rect 5458 21758 5460 21810
rect 5404 21746 5460 21758
rect 4676 21532 4900 21588
rect 4620 21494 4676 21532
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 3612 20802 3668 20814
rect 3612 20750 3614 20802
rect 3666 20750 3668 20802
rect 3612 20580 3668 20750
rect 4732 20692 4788 20702
rect 3612 20514 3668 20524
rect 3836 20580 3892 20590
rect 4172 20580 4228 20590
rect 3836 20578 4004 20580
rect 3836 20526 3838 20578
rect 3890 20526 4004 20578
rect 3836 20524 4004 20526
rect 3836 20514 3892 20524
rect 3276 20412 3444 20468
rect 3164 19460 3220 20188
rect 3276 20132 3332 20142
rect 3276 20038 3332 20076
rect 3276 19460 3332 19470
rect 3164 19458 3332 19460
rect 3164 19406 3278 19458
rect 3330 19406 3332 19458
rect 3164 19404 3332 19406
rect 3276 19394 3332 19404
rect 3052 19348 3108 19358
rect 2940 19346 3108 19348
rect 2940 19294 3054 19346
rect 3106 19294 3108 19346
rect 2940 19292 3108 19294
rect 2044 19124 2100 19134
rect 2940 19124 2996 19292
rect 3052 19282 3108 19292
rect 3388 19236 3444 20412
rect 3836 20244 3892 20254
rect 3836 20150 3892 20188
rect 3724 20132 3780 20142
rect 3724 20038 3780 20076
rect 3948 20020 4004 20524
rect 4060 20020 4116 20030
rect 3948 19964 4060 20020
rect 4060 19954 4116 19964
rect 2044 19122 2996 19124
rect 2044 19070 2046 19122
rect 2098 19070 2996 19122
rect 2044 19068 2996 19070
rect 3164 19180 3444 19236
rect 4172 19234 4228 20524
rect 4508 20580 4564 20590
rect 4508 20486 4564 20524
rect 4172 19182 4174 19234
rect 4226 19182 4228 19234
rect 2044 19058 2100 19068
rect 1932 18386 1988 18396
rect 3164 16884 3220 19180
rect 4172 19170 4228 19182
rect 4284 20018 4340 20030
rect 4284 19966 4286 20018
rect 4338 19966 4340 20018
rect 3612 19012 3668 19022
rect 3612 18918 3668 18956
rect 4284 18900 4340 19966
rect 4732 20018 4788 20636
rect 4844 20356 4900 21532
rect 5180 21586 5348 21588
rect 5180 21534 5182 21586
rect 5234 21534 5348 21586
rect 5180 21532 5348 21534
rect 4956 21028 5012 21038
rect 5180 21028 5236 21532
rect 5516 21474 5572 22652
rect 5628 21586 5684 22764
rect 5740 21812 5796 23102
rect 5740 21746 5796 21756
rect 5628 21534 5630 21586
rect 5682 21534 5684 21586
rect 5628 21522 5684 21534
rect 5852 21700 5908 21710
rect 5516 21422 5518 21474
rect 5570 21422 5572 21474
rect 5516 21410 5572 21422
rect 5740 21028 5796 21038
rect 5180 21026 5796 21028
rect 5180 20974 5742 21026
rect 5794 20974 5796 21026
rect 5180 20972 5796 20974
rect 4956 20934 5012 20972
rect 5740 20962 5796 20972
rect 5852 21026 5908 21644
rect 5852 20974 5854 21026
rect 5906 20974 5908 21026
rect 5852 20962 5908 20974
rect 5964 21586 6020 23214
rect 6412 23156 6468 23774
rect 6524 23716 6580 23726
rect 6524 23622 6580 23660
rect 6524 23380 6580 23390
rect 6636 23380 6692 23884
rect 6748 23938 6804 23996
rect 6748 23886 6750 23938
rect 6802 23886 6804 23938
rect 6748 23874 6804 23886
rect 7420 23492 7476 24670
rect 7644 24722 7700 24734
rect 7644 24670 7646 24722
rect 7698 24670 7700 24722
rect 7532 24612 7588 24622
rect 7532 24518 7588 24556
rect 7420 23426 7476 23436
rect 6524 23378 6692 23380
rect 6524 23326 6526 23378
rect 6578 23326 6692 23378
rect 6524 23324 6692 23326
rect 6524 23314 6580 23324
rect 6412 23100 6580 23156
rect 6412 22930 6468 22942
rect 6412 22878 6414 22930
rect 6466 22878 6468 22930
rect 6412 22820 6468 22878
rect 6412 22754 6468 22764
rect 6524 22708 6580 23100
rect 6524 22642 6580 22652
rect 6636 22932 6692 23324
rect 7196 23380 7252 23390
rect 7196 23286 7252 23324
rect 7644 23380 7700 24670
rect 7644 23314 7700 23324
rect 7756 24722 7812 24734
rect 7756 24670 7758 24722
rect 7810 24670 7812 24722
rect 7756 23714 7812 24670
rect 8652 24722 8708 25228
rect 9212 25284 9268 25294
rect 9212 25190 9268 25228
rect 8652 24670 8654 24722
rect 8706 24670 8708 24722
rect 8652 24658 8708 24670
rect 8652 24498 8708 24510
rect 8652 24446 8654 24498
rect 8706 24446 8708 24498
rect 8540 24050 8596 24062
rect 8540 23998 8542 24050
rect 8594 23998 8596 24050
rect 7980 23940 8036 23950
rect 7980 23846 8036 23884
rect 7756 23662 7758 23714
rect 7810 23662 7812 23714
rect 7420 23268 7476 23278
rect 7420 23174 7476 23212
rect 7084 23154 7140 23166
rect 7084 23102 7086 23154
rect 7138 23102 7140 23154
rect 6412 22596 6468 22606
rect 6300 22484 6356 22494
rect 6300 22370 6356 22428
rect 6412 22482 6468 22540
rect 6412 22430 6414 22482
rect 6466 22430 6468 22482
rect 6412 22418 6468 22430
rect 6636 22484 6692 22876
rect 6636 22418 6692 22428
rect 6748 22930 6804 22942
rect 6748 22878 6750 22930
rect 6802 22878 6804 22930
rect 6300 22318 6302 22370
rect 6354 22318 6356 22370
rect 6300 22306 6356 22318
rect 6748 22372 6804 22878
rect 6748 22306 6804 22316
rect 5964 21534 5966 21586
rect 6018 21534 6020 21586
rect 5068 20690 5124 20702
rect 5964 20692 6020 21534
rect 6188 22258 6244 22270
rect 6188 22206 6190 22258
rect 6242 22206 6244 22258
rect 6188 21586 6244 22206
rect 6524 22148 6580 22158
rect 6524 22054 6580 22092
rect 6748 22148 6804 22158
rect 6748 22146 6916 22148
rect 6748 22094 6750 22146
rect 6802 22094 6916 22146
rect 6748 22092 6916 22094
rect 6748 22082 6804 22092
rect 6748 21924 6804 21934
rect 6748 21810 6804 21868
rect 6748 21758 6750 21810
rect 6802 21758 6804 21810
rect 6748 21746 6804 21758
rect 6860 21810 6916 22092
rect 7084 21924 7140 23102
rect 7084 21858 7140 21868
rect 6860 21758 6862 21810
rect 6914 21758 6916 21810
rect 6636 21700 6692 21710
rect 6636 21606 6692 21644
rect 6188 21534 6190 21586
rect 6242 21534 6244 21586
rect 6188 21028 6244 21534
rect 6188 20962 6244 20972
rect 6748 21476 6804 21486
rect 6076 20804 6132 20814
rect 6076 20710 6132 20748
rect 6188 20802 6244 20814
rect 6188 20750 6190 20802
rect 6242 20750 6244 20802
rect 5068 20638 5070 20690
rect 5122 20638 5124 20690
rect 4844 20290 4900 20300
rect 4956 20578 5012 20590
rect 4956 20526 4958 20578
rect 5010 20526 5012 20578
rect 4732 19966 4734 20018
rect 4786 19966 4788 20018
rect 4732 19908 4788 19966
rect 4956 20020 5012 20526
rect 5068 20356 5124 20638
rect 5740 20636 6020 20692
rect 5068 20300 5684 20356
rect 4956 19954 5012 19964
rect 4732 19842 4788 19852
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4620 19460 4676 19470
rect 4620 19234 4676 19404
rect 4732 19348 4788 19358
rect 4732 19254 4788 19292
rect 4620 19182 4622 19234
rect 4674 19182 4676 19234
rect 4620 19170 4676 19182
rect 4284 18844 4452 18900
rect 3836 18676 3892 18686
rect 4284 18676 4340 18686
rect 3836 18674 4340 18676
rect 3836 18622 3838 18674
rect 3890 18622 4286 18674
rect 4338 18622 4340 18674
rect 3836 18620 4340 18622
rect 3836 18610 3892 18620
rect 4284 18610 4340 18620
rect 3724 18452 3780 18462
rect 3724 18358 3780 18396
rect 4172 18452 4228 18462
rect 4172 18358 4228 18396
rect 4396 18228 4452 18844
rect 5180 18674 5236 20300
rect 5628 20242 5684 20300
rect 5628 20190 5630 20242
rect 5682 20190 5684 20242
rect 5628 20178 5684 20190
rect 5740 20242 5796 20636
rect 5740 20190 5742 20242
rect 5794 20190 5796 20242
rect 5740 20178 5796 20190
rect 5852 20468 5908 20478
rect 5292 20132 5348 20142
rect 5348 20076 5460 20132
rect 5292 20038 5348 20076
rect 5180 18622 5182 18674
rect 5234 18622 5236 18674
rect 5180 18610 5236 18622
rect 5292 19908 5348 19918
rect 5292 18674 5348 19852
rect 5404 19236 5460 20076
rect 5852 20018 5908 20412
rect 6188 20244 6244 20750
rect 6636 20804 6692 20814
rect 6636 20710 6692 20748
rect 6748 20692 6804 21420
rect 6860 20914 6916 21758
rect 7196 21812 7252 21822
rect 7196 21476 7252 21756
rect 7532 21700 7588 21710
rect 7532 21606 7588 21644
rect 7196 21410 7252 21420
rect 6860 20862 6862 20914
rect 6914 20862 6916 20914
rect 6860 20850 6916 20862
rect 6972 20692 7028 20702
rect 6748 20636 6916 20692
rect 5852 19966 5854 20018
rect 5906 19966 5908 20018
rect 5740 19460 5796 19470
rect 5852 19460 5908 19966
rect 5740 19458 5908 19460
rect 5740 19406 5742 19458
rect 5794 19406 5908 19458
rect 5740 19404 5908 19406
rect 5964 20188 6244 20244
rect 6860 20242 6916 20636
rect 6972 20690 7700 20692
rect 6972 20638 6974 20690
rect 7026 20638 7700 20690
rect 6972 20636 7700 20638
rect 6972 20626 7028 20636
rect 6860 20190 6862 20242
rect 6914 20190 6916 20242
rect 5740 19394 5796 19404
rect 5628 19236 5684 19246
rect 5404 19234 5684 19236
rect 5404 19182 5630 19234
rect 5682 19182 5684 19234
rect 5404 19180 5684 19182
rect 5628 19170 5684 19180
rect 5292 18622 5294 18674
rect 5346 18622 5348 18674
rect 5292 18610 5348 18622
rect 5404 18788 5460 18798
rect 4172 18172 4452 18228
rect 4508 18450 4564 18462
rect 4508 18398 4510 18450
rect 4562 18398 4564 18450
rect 4508 18228 4564 18398
rect 4172 17332 4228 18172
rect 4508 18162 4564 18172
rect 5404 18228 5460 18732
rect 5516 18452 5572 18462
rect 5516 18450 5684 18452
rect 5516 18398 5518 18450
rect 5570 18398 5684 18450
rect 5516 18396 5684 18398
rect 5516 18386 5572 18396
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4172 17276 4452 17332
rect 3276 16884 3332 16894
rect 3164 16882 3332 16884
rect 3164 16830 3278 16882
rect 3330 16830 3332 16882
rect 3164 16828 3332 16830
rect 3276 16818 3332 16828
rect 3276 16660 3332 16670
rect 2492 16658 3332 16660
rect 2492 16606 3278 16658
rect 3330 16606 3332 16658
rect 2492 16604 3332 16606
rect 2492 16210 2548 16604
rect 3276 16594 3332 16604
rect 3612 16660 3668 16670
rect 3612 16566 3668 16604
rect 4284 16324 4340 17276
rect 4396 17106 4452 17276
rect 4396 17054 4398 17106
rect 4450 17054 4452 17106
rect 4396 17042 4452 17054
rect 4732 16994 4788 17006
rect 4732 16942 4734 16994
rect 4786 16942 4788 16994
rect 4732 16660 4788 16942
rect 4732 16604 4900 16660
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4844 16436 4900 16604
rect 4844 16370 4900 16380
rect 4956 16548 5012 16558
rect 4620 16324 4676 16334
rect 4284 16268 4620 16324
rect 2492 16158 2494 16210
rect 2546 16158 2548 16210
rect 2492 16146 2548 16158
rect 4620 16210 4676 16268
rect 4620 16158 4622 16210
rect 4674 16158 4676 16210
rect 4620 16146 4676 16158
rect 1820 16098 1876 16110
rect 1820 16046 1822 16098
rect 1874 16046 1876 16098
rect 1820 13746 1876 16046
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4956 14642 5012 16492
rect 5068 15876 5124 15886
rect 5068 15874 5348 15876
rect 5068 15822 5070 15874
rect 5122 15822 5348 15874
rect 5068 15820 5348 15822
rect 5068 15810 5124 15820
rect 4956 14590 4958 14642
rect 5010 14590 5012 14642
rect 4956 14578 5012 14590
rect 5068 14644 5124 14682
rect 5068 14578 5124 14588
rect 4844 14532 4900 14542
rect 4844 14418 4900 14476
rect 4844 14366 4846 14418
rect 4898 14366 4900 14418
rect 4844 14354 4900 14366
rect 5292 14084 5348 15820
rect 5404 15540 5460 18172
rect 5628 17444 5684 18396
rect 5852 18450 5908 18462
rect 5852 18398 5854 18450
rect 5906 18398 5908 18450
rect 5628 17388 5796 17444
rect 5628 17220 5684 17230
rect 5516 17164 5628 17220
rect 5516 16322 5572 17164
rect 5628 17154 5684 17164
rect 5740 16994 5796 17388
rect 5740 16942 5742 16994
rect 5794 16942 5796 16994
rect 5628 16882 5684 16894
rect 5628 16830 5630 16882
rect 5682 16830 5684 16882
rect 5628 16548 5684 16830
rect 5628 16482 5684 16492
rect 5740 16436 5796 16942
rect 5852 16548 5908 18398
rect 5964 17666 6020 20188
rect 6860 20178 6916 20190
rect 6636 20130 6692 20142
rect 6636 20078 6638 20130
rect 6690 20078 6692 20130
rect 6188 20020 6244 20030
rect 6076 18900 6132 18910
rect 6076 18562 6132 18844
rect 6076 18510 6078 18562
rect 6130 18510 6132 18562
rect 6076 18498 6132 18510
rect 6188 18340 6244 19964
rect 6524 20018 6580 20030
rect 6524 19966 6526 20018
rect 6578 19966 6580 20018
rect 6524 19460 6580 19966
rect 6524 19394 6580 19404
rect 6636 19236 6692 20078
rect 6524 19180 6692 19236
rect 7644 19236 7700 20636
rect 7756 19908 7812 23662
rect 8428 22372 8484 22382
rect 8428 20242 8484 22316
rect 8540 20692 8596 23998
rect 8652 23940 8708 24446
rect 8652 23874 8708 23884
rect 8988 24498 9044 24510
rect 8988 24446 8990 24498
rect 9042 24446 9044 24498
rect 8876 23604 8932 23614
rect 8876 23266 8932 23548
rect 8876 23214 8878 23266
rect 8930 23214 8932 23266
rect 8652 22930 8708 22942
rect 8652 22878 8654 22930
rect 8706 22878 8708 22930
rect 8652 22372 8708 22878
rect 8652 22306 8708 22316
rect 8876 20916 8932 23214
rect 8988 22932 9044 24446
rect 8988 22930 9156 22932
rect 8988 22878 8990 22930
rect 9042 22878 9156 22930
rect 8988 22876 9156 22878
rect 8988 22866 9044 22876
rect 8988 20916 9044 20926
rect 8876 20860 8988 20916
rect 8988 20850 9044 20860
rect 8540 20626 8596 20636
rect 8428 20190 8430 20242
rect 8482 20190 8484 20242
rect 8428 20178 8484 20190
rect 8204 20020 8260 20030
rect 8540 20020 8596 20030
rect 8204 19926 8260 19964
rect 8428 20018 8596 20020
rect 8428 19966 8542 20018
rect 8594 19966 8596 20018
rect 8428 19964 8596 19966
rect 8428 19908 8484 19964
rect 8540 19954 8596 19964
rect 8652 20020 8708 20030
rect 8652 19926 8708 19964
rect 8988 20018 9044 20030
rect 8988 19966 8990 20018
rect 9042 19966 9044 20018
rect 7756 19852 8036 19908
rect 7868 19236 7924 19246
rect 7644 19234 7924 19236
rect 7644 19182 7870 19234
rect 7922 19182 7924 19234
rect 7644 19180 7924 19182
rect 6300 19122 6356 19134
rect 6300 19070 6302 19122
rect 6354 19070 6356 19122
rect 6300 19012 6356 19070
rect 6300 18946 6356 18956
rect 6412 19124 6468 19134
rect 6524 19124 6580 19180
rect 6468 19068 6580 19124
rect 7308 19122 7364 19134
rect 7308 19070 7310 19122
rect 7362 19070 7364 19122
rect 6412 19010 6468 19068
rect 6412 18958 6414 19010
rect 6466 18958 6468 19010
rect 6412 18788 6468 18958
rect 6636 19012 6692 19022
rect 6636 18918 6692 18956
rect 6412 18722 6468 18732
rect 6300 18564 6356 18574
rect 6300 18470 6356 18508
rect 7196 18452 7252 18462
rect 7084 18396 7196 18452
rect 6188 18284 6356 18340
rect 5964 17614 5966 17666
rect 6018 17614 6020 17666
rect 5964 17220 6020 17614
rect 6188 18004 6244 18014
rect 6188 17554 6244 17948
rect 6188 17502 6190 17554
rect 6242 17502 6244 17554
rect 6188 17490 6244 17502
rect 5964 17154 6020 17164
rect 6300 16994 6356 18284
rect 6412 18228 6468 18238
rect 6412 18226 7028 18228
rect 6412 18174 6414 18226
rect 6466 18174 7028 18226
rect 6412 18172 7028 18174
rect 6412 18162 6468 18172
rect 6860 18004 6916 18014
rect 6860 17666 6916 17948
rect 6860 17614 6862 17666
rect 6914 17614 6916 17666
rect 6860 17602 6916 17614
rect 6972 17554 7028 18172
rect 6972 17502 6974 17554
rect 7026 17502 7028 17554
rect 6972 17490 7028 17502
rect 6524 17108 6580 17118
rect 7084 17108 7140 18396
rect 7196 18358 7252 18396
rect 7308 18338 7364 19070
rect 7532 19124 7588 19134
rect 7532 19030 7588 19068
rect 7420 19012 7476 19022
rect 7420 18674 7476 18956
rect 7644 18788 7700 19180
rect 7868 19170 7924 19180
rect 7756 19012 7812 19022
rect 7756 18918 7812 18956
rect 7420 18622 7422 18674
rect 7474 18622 7476 18674
rect 7420 18610 7476 18622
rect 7532 18732 7700 18788
rect 7308 18286 7310 18338
rect 7362 18286 7364 18338
rect 7308 18274 7364 18286
rect 7532 18228 7588 18732
rect 7644 18564 7700 18574
rect 7644 18470 7700 18508
rect 7868 18452 7924 18462
rect 7532 18162 7588 18172
rect 7756 18450 7924 18452
rect 7756 18398 7870 18450
rect 7922 18398 7924 18450
rect 7756 18396 7924 18398
rect 7756 18004 7812 18396
rect 7868 18386 7924 18396
rect 7196 17948 7812 18004
rect 7196 17666 7252 17948
rect 7196 17614 7198 17666
rect 7250 17614 7252 17666
rect 7196 17602 7252 17614
rect 6524 17106 7140 17108
rect 6524 17054 6526 17106
rect 6578 17054 7140 17106
rect 6524 17052 7140 17054
rect 6524 17042 6580 17052
rect 6300 16942 6302 16994
rect 6354 16942 6356 16994
rect 5964 16884 6020 16894
rect 6188 16884 6244 16894
rect 5964 16882 6244 16884
rect 5964 16830 5966 16882
rect 6018 16830 6190 16882
rect 6242 16830 6244 16882
rect 5964 16828 6244 16830
rect 5964 16818 6020 16828
rect 6188 16818 6244 16828
rect 5852 16482 5908 16492
rect 5740 16370 5796 16380
rect 5516 16270 5518 16322
rect 5570 16270 5572 16322
rect 5516 16258 5572 16270
rect 6188 16324 6244 16334
rect 6188 16230 6244 16268
rect 5964 16098 6020 16110
rect 5964 16046 5966 16098
rect 6018 16046 6020 16098
rect 5628 15540 5684 15550
rect 5404 15538 5684 15540
rect 5404 15486 5630 15538
rect 5682 15486 5684 15538
rect 5404 15484 5684 15486
rect 5628 15474 5684 15484
rect 5964 15540 6020 16046
rect 5964 15474 6020 15484
rect 6188 15540 6244 15550
rect 6300 15540 6356 16942
rect 7084 16884 7140 17052
rect 7308 16884 7364 16894
rect 7532 16884 7588 16922
rect 7084 16882 7364 16884
rect 7084 16830 7310 16882
rect 7362 16830 7364 16882
rect 7084 16828 7364 16830
rect 7308 16818 7364 16828
rect 7420 16828 7532 16884
rect 7084 16658 7140 16670
rect 7084 16606 7086 16658
rect 7138 16606 7140 16658
rect 6748 16548 6804 16558
rect 6748 16322 6804 16492
rect 6748 16270 6750 16322
rect 6802 16270 6804 16322
rect 6748 16258 6804 16270
rect 7084 16322 7140 16606
rect 7084 16270 7086 16322
rect 7138 16270 7140 16322
rect 7084 16258 7140 16270
rect 7308 16212 7364 16222
rect 6412 16100 6468 16110
rect 6412 16006 6468 16044
rect 7084 16100 7140 16110
rect 6188 15538 6356 15540
rect 6188 15486 6190 15538
rect 6242 15486 6356 15538
rect 6188 15484 6356 15486
rect 6972 15988 7028 15998
rect 6972 15874 7028 15932
rect 6972 15822 6974 15874
rect 7026 15822 7028 15874
rect 6188 15474 6244 15484
rect 5516 15316 5572 15326
rect 5516 15222 5572 15260
rect 6076 15314 6132 15326
rect 6076 15262 6078 15314
rect 6130 15262 6132 15314
rect 5628 15092 5684 15102
rect 5628 15090 5796 15092
rect 5628 15038 5630 15090
rect 5682 15038 5796 15090
rect 5628 15036 5796 15038
rect 5628 15026 5684 15036
rect 5068 14028 5348 14084
rect 5516 14644 5572 14654
rect 5068 13972 5124 14028
rect 4956 13970 5124 13972
rect 4956 13918 5070 13970
rect 5122 13918 5124 13970
rect 4956 13916 5124 13918
rect 2492 13860 2548 13870
rect 2492 13766 2548 13804
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 11396 1876 13694
rect 4620 13636 4676 13646
rect 4620 13634 4900 13636
rect 4620 13582 4622 13634
rect 4674 13582 4900 13634
rect 4620 13580 4900 13582
rect 4620 13570 4676 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4844 12964 4900 13580
rect 4844 12898 4900 12908
rect 4844 12292 4900 12302
rect 4844 12178 4900 12236
rect 4844 12126 4846 12178
rect 4898 12126 4900 12178
rect 4508 12068 4564 12078
rect 4508 11974 4564 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11506 4900 12126
rect 4844 11454 4846 11506
rect 4898 11454 4900 11506
rect 4844 11442 4900 11454
rect 4956 12068 5012 13916
rect 5068 13906 5124 13916
rect 5516 13188 5572 14588
rect 5740 13858 5796 15036
rect 6076 14756 6132 15262
rect 6972 15204 7028 15822
rect 6972 15138 7028 15148
rect 7084 15428 7140 16044
rect 6188 15092 6244 15102
rect 6188 15090 6356 15092
rect 6188 15038 6190 15090
rect 6242 15038 6356 15090
rect 6188 15036 6356 15038
rect 6188 15026 6244 15036
rect 5852 14700 6132 14756
rect 5852 14644 5908 14700
rect 6188 14644 6244 14654
rect 5852 14578 5908 14588
rect 6076 14642 6244 14644
rect 6076 14590 6190 14642
rect 6242 14590 6244 14642
rect 6076 14588 6244 14590
rect 5964 14532 6020 14542
rect 5964 14438 6020 14476
rect 6076 13970 6132 14588
rect 6188 14578 6244 14588
rect 6076 13918 6078 13970
rect 6130 13918 6132 13970
rect 6076 13906 6132 13918
rect 5740 13806 5742 13858
rect 5794 13806 5796 13858
rect 5740 13794 5796 13806
rect 5852 13858 5908 13870
rect 5852 13806 5854 13858
rect 5906 13806 5908 13858
rect 5740 13188 5796 13198
rect 5516 13186 5796 13188
rect 5516 13134 5742 13186
rect 5794 13134 5796 13186
rect 5516 13132 5796 13134
rect 5740 13122 5796 13132
rect 5852 13076 5908 13806
rect 5852 13010 5908 13020
rect 6188 13076 6244 13086
rect 6300 13076 6356 15036
rect 7084 14642 7140 15372
rect 7196 15314 7252 15326
rect 7196 15262 7198 15314
rect 7250 15262 7252 15314
rect 7196 15204 7252 15262
rect 7196 15138 7252 15148
rect 7084 14590 7086 14642
rect 7138 14590 7140 14642
rect 7084 14578 7140 14590
rect 6972 14532 7028 14542
rect 6972 14438 7028 14476
rect 6636 14420 6692 14430
rect 6636 14326 6692 14364
rect 6244 13020 6356 13076
rect 6188 13010 6244 13020
rect 5516 12964 5572 12974
rect 5292 12908 5516 12964
rect 5292 12180 5348 12908
rect 5516 12870 5572 12908
rect 5852 12738 5908 12750
rect 5852 12686 5854 12738
rect 5906 12686 5908 12738
rect 5740 12180 5796 12190
rect 5292 12178 5684 12180
rect 5292 12126 5294 12178
rect 5346 12126 5684 12178
rect 5292 12124 5684 12126
rect 5292 12114 5348 12124
rect 2044 11396 2100 11406
rect 1820 11394 2100 11396
rect 1820 11342 2046 11394
rect 2098 11342 2100 11394
rect 1820 11340 2100 11342
rect 2044 10612 2100 11340
rect 2716 11282 2772 11294
rect 2716 11230 2718 11282
rect 2770 11230 2772 11282
rect 2716 10836 2772 11230
rect 2716 10770 2772 10780
rect 4956 10836 5012 12012
rect 2380 10612 2436 10622
rect 2044 10610 2436 10612
rect 2044 10558 2382 10610
rect 2434 10558 2436 10610
rect 2044 10556 2436 10558
rect 2380 10500 2436 10556
rect 3052 10612 3108 10622
rect 3052 10518 3108 10556
rect 2380 10434 2436 10444
rect 4956 10500 5012 10780
rect 5068 11954 5124 11966
rect 5068 11902 5070 11954
rect 5122 11902 5124 11954
rect 5068 10500 5124 11902
rect 5628 11394 5684 12124
rect 5740 12086 5796 12124
rect 5628 11342 5630 11394
rect 5682 11342 5684 11394
rect 5628 11330 5684 11342
rect 5852 11732 5908 12686
rect 6076 12738 6132 12750
rect 6076 12686 6078 12738
rect 6130 12686 6132 12738
rect 6076 12516 6132 12686
rect 6076 12460 6356 12516
rect 6076 12292 6132 12460
rect 6300 12402 6356 12460
rect 6300 12350 6302 12402
rect 6354 12350 6356 12402
rect 6300 12338 6356 12350
rect 6636 12404 6692 12414
rect 6636 12310 6692 12348
rect 6076 12226 6132 12236
rect 5852 10834 5908 11676
rect 6748 11956 6804 11966
rect 6748 11394 6804 11900
rect 6748 11342 6750 11394
rect 6802 11342 6804 11394
rect 5964 11284 6020 11294
rect 5964 11190 6020 11228
rect 6748 11284 6804 11342
rect 7196 11732 7252 11742
rect 7196 11394 7252 11676
rect 7196 11342 7198 11394
rect 7250 11342 7252 11394
rect 7196 11330 7252 11342
rect 6748 11218 6804 11228
rect 5852 10782 5854 10834
rect 5906 10782 5908 10834
rect 5852 10770 5908 10782
rect 6300 10836 6356 10846
rect 5516 10610 5572 10622
rect 5516 10558 5518 10610
rect 5570 10558 5572 10610
rect 5180 10500 5236 10510
rect 5516 10500 5572 10558
rect 5068 10498 5572 10500
rect 5068 10446 5182 10498
rect 5234 10446 5572 10498
rect 5068 10444 5572 10446
rect 4956 10434 5012 10444
rect 5180 10434 5236 10444
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 6300 8372 6356 10780
rect 7308 10610 7364 16156
rect 7420 13860 7476 16828
rect 7532 16818 7588 16828
rect 7756 16884 7812 16894
rect 7756 16790 7812 16828
rect 7644 16770 7700 16782
rect 7644 16718 7646 16770
rect 7698 16718 7700 16770
rect 7532 16660 7588 16670
rect 7532 16210 7588 16604
rect 7644 16324 7700 16718
rect 7644 16268 7924 16324
rect 7532 16158 7534 16210
rect 7586 16158 7588 16210
rect 7532 16146 7588 16158
rect 7868 16098 7924 16268
rect 7868 16046 7870 16098
rect 7922 16046 7924 16098
rect 7868 16034 7924 16046
rect 7644 15988 7700 15998
rect 7644 15894 7700 15932
rect 7532 15874 7588 15886
rect 7532 15822 7534 15874
rect 7586 15822 7588 15874
rect 7532 15764 7588 15822
rect 7980 15764 8036 19852
rect 8428 19842 8484 19852
rect 8988 19908 9044 19966
rect 8988 19842 9044 19852
rect 8316 19236 8372 19246
rect 8316 19142 8372 19180
rect 8988 19236 9044 19246
rect 8988 19142 9044 19180
rect 8204 19010 8260 19022
rect 8204 18958 8206 19010
rect 8258 18958 8260 19010
rect 8204 18674 8260 18958
rect 8428 19012 8484 19022
rect 8428 18918 8484 18956
rect 8652 19010 8708 19022
rect 8652 18958 8654 19010
rect 8706 18958 8708 19010
rect 8652 18900 8708 18958
rect 8652 18834 8708 18844
rect 8988 18900 9044 18910
rect 8204 18622 8206 18674
rect 8258 18622 8260 18674
rect 8204 18610 8260 18622
rect 8988 18674 9044 18844
rect 8988 18622 8990 18674
rect 9042 18622 9044 18674
rect 8988 18610 9044 18622
rect 8428 18564 8484 18574
rect 8204 18452 8260 18462
rect 8204 18358 8260 18396
rect 8428 18450 8484 18508
rect 8428 18398 8430 18450
rect 8482 18398 8484 18450
rect 8428 18386 8484 18398
rect 8204 18228 8260 18238
rect 8204 16882 8260 18172
rect 8204 16830 8206 16882
rect 8258 16830 8260 16882
rect 8204 16818 8260 16830
rect 8764 16884 8820 16894
rect 8764 16790 8820 16828
rect 8428 16660 8484 16670
rect 8316 16658 8484 16660
rect 8316 16606 8430 16658
rect 8482 16606 8484 16658
rect 8316 16604 8484 16606
rect 8092 16212 8148 16222
rect 8092 16098 8148 16156
rect 8092 16046 8094 16098
rect 8146 16046 8148 16098
rect 8092 16034 8148 16046
rect 7532 15708 8148 15764
rect 7756 15540 7812 15550
rect 7756 15446 7812 15484
rect 7644 15428 7700 15438
rect 7644 15334 7700 15372
rect 7868 15316 7924 15354
rect 7756 15260 7868 15316
rect 7532 13860 7588 13870
rect 7420 13858 7588 13860
rect 7420 13806 7534 13858
rect 7586 13806 7588 13858
rect 7420 13804 7588 13806
rect 7532 13794 7588 13804
rect 7420 13188 7476 13198
rect 7420 13094 7476 13132
rect 7644 13076 7700 13086
rect 7644 12982 7700 13020
rect 7756 12180 7812 15260
rect 7868 15250 7924 15260
rect 8092 13970 8148 15708
rect 8316 15540 8372 16604
rect 8428 16594 8484 16604
rect 9100 16548 9156 22876
rect 9212 20692 9268 20702
rect 9212 19684 9268 20636
rect 9436 20580 9492 27356
rect 10332 27298 10388 27804
rect 10556 27636 10612 30268
rect 10892 30258 10948 30268
rect 10780 29314 10836 29326
rect 10780 29262 10782 29314
rect 10834 29262 10836 29314
rect 10780 29204 10836 29262
rect 11004 29204 11060 30940
rect 11452 30930 11508 30940
rect 10836 29148 11060 29204
rect 11116 29428 11172 29438
rect 10780 29110 10836 29148
rect 11116 28868 11172 29372
rect 11564 29204 11620 32956
rect 11676 32946 11732 32956
rect 12236 33236 12292 33246
rect 12236 32450 12292 33180
rect 12236 32398 12238 32450
rect 12290 32398 12292 32450
rect 11676 32004 11732 32014
rect 11676 31218 11732 31948
rect 11676 31166 11678 31218
rect 11730 31166 11732 31218
rect 11676 31154 11732 31166
rect 12236 30994 12292 32398
rect 12796 31890 12852 34860
rect 13244 34354 13300 34860
rect 13244 34302 13246 34354
rect 13298 34302 13300 34354
rect 13244 34290 13300 34302
rect 13580 34692 13636 34702
rect 13580 34354 13636 34636
rect 13580 34302 13582 34354
rect 13634 34302 13636 34354
rect 13580 34290 13636 34302
rect 13468 33460 13524 33470
rect 12796 31838 12798 31890
rect 12850 31838 12852 31890
rect 12796 31826 12852 31838
rect 12908 33458 13524 33460
rect 12908 33406 13470 33458
rect 13522 33406 13524 33458
rect 12908 33404 13524 33406
rect 12684 31668 12740 31678
rect 12684 31574 12740 31612
rect 12908 31106 12964 33404
rect 13468 33394 13524 33404
rect 13580 33236 13636 33246
rect 13692 33236 13748 35420
rect 14028 35382 14084 35420
rect 14588 34916 14644 36206
rect 14700 34916 14756 34926
rect 14588 34914 14756 34916
rect 14588 34862 14702 34914
rect 14754 34862 14756 34914
rect 14588 34860 14756 34862
rect 14700 34850 14756 34860
rect 14812 34692 14868 36876
rect 14924 36706 14980 37100
rect 14924 36654 14926 36706
rect 14978 36654 14980 36706
rect 14924 36642 14980 36654
rect 15036 36148 15092 37548
rect 15260 37492 15316 37884
rect 15484 37874 15540 37884
rect 15148 36596 15204 36606
rect 15260 36596 15316 37436
rect 15596 37826 15652 37838
rect 15596 37774 15598 37826
rect 15650 37774 15652 37826
rect 15484 37268 15540 37278
rect 15484 37174 15540 37212
rect 15596 37044 15652 37774
rect 15820 37828 15876 37838
rect 15820 37734 15876 37772
rect 16268 37492 16324 38110
rect 21532 38164 21588 38174
rect 21532 38162 21812 38164
rect 21532 38110 21534 38162
rect 21586 38110 21812 38162
rect 21532 38108 21812 38110
rect 21532 38098 21588 38108
rect 19180 38050 19236 38062
rect 19180 37998 19182 38050
rect 19234 37998 19236 38050
rect 18396 37940 18452 37950
rect 17724 37938 18452 37940
rect 17724 37886 18398 37938
rect 18450 37886 18452 37938
rect 17724 37884 18452 37886
rect 16044 37436 16324 37492
rect 16716 37828 16772 37838
rect 15708 37154 15764 37166
rect 15708 37102 15710 37154
rect 15762 37102 15764 37154
rect 15708 37044 15764 37102
rect 16044 37044 16100 37436
rect 16716 37378 16772 37772
rect 17612 37828 17668 37838
rect 17612 37490 17668 37772
rect 17612 37438 17614 37490
rect 17666 37438 17668 37490
rect 17612 37426 17668 37438
rect 16716 37326 16718 37378
rect 16770 37326 16772 37378
rect 16716 37314 16772 37326
rect 17388 37378 17444 37390
rect 17388 37326 17390 37378
rect 17442 37326 17444 37378
rect 16156 37266 16212 37278
rect 16380 37268 16436 37278
rect 16156 37214 16158 37266
rect 16210 37214 16212 37266
rect 16156 37156 16212 37214
rect 16156 37090 16212 37100
rect 16268 37212 16380 37268
rect 15708 36988 16100 37044
rect 15596 36978 15652 36988
rect 15148 36594 15316 36596
rect 15148 36542 15150 36594
rect 15202 36542 15316 36594
rect 15148 36540 15316 36542
rect 15148 36530 15204 36540
rect 15484 36484 15540 36494
rect 15932 36484 15988 36988
rect 16044 36484 16100 36494
rect 15932 36428 16044 36484
rect 15148 36148 15204 36158
rect 15036 36092 15148 36148
rect 15148 36082 15204 36092
rect 15260 35028 15316 35038
rect 15260 35026 15428 35028
rect 15260 34974 15262 35026
rect 15314 34974 15428 35026
rect 15260 34972 15428 34974
rect 15260 34962 15316 34972
rect 14924 34692 14980 34702
rect 14812 34690 14980 34692
rect 14812 34638 14926 34690
rect 14978 34638 14980 34690
rect 14812 34636 14980 34638
rect 14924 34580 14980 34636
rect 15148 34692 15204 34702
rect 15148 34598 15204 34636
rect 15260 34690 15316 34702
rect 15260 34638 15262 34690
rect 15314 34638 15316 34690
rect 14924 34514 14980 34524
rect 15260 34468 15316 34638
rect 15260 34402 15316 34412
rect 14924 34244 14980 34254
rect 15372 34244 15428 34972
rect 13804 34020 13860 34030
rect 13804 33570 13860 33964
rect 13804 33518 13806 33570
rect 13858 33518 13860 33570
rect 13804 33506 13860 33518
rect 14252 34018 14308 34030
rect 14252 33966 14254 34018
rect 14306 33966 14308 34018
rect 13580 33234 13748 33236
rect 13580 33182 13582 33234
rect 13634 33182 13748 33234
rect 13580 33180 13748 33182
rect 14252 33236 14308 33966
rect 14812 33460 14868 33470
rect 14812 33346 14868 33404
rect 14924 33458 14980 34188
rect 14924 33406 14926 33458
rect 14978 33406 14980 33458
rect 14924 33394 14980 33406
rect 15036 34188 15428 34244
rect 14812 33294 14814 33346
rect 14866 33294 14868 33346
rect 14812 33282 14868 33294
rect 15036 33346 15092 34188
rect 15372 34130 15428 34188
rect 15372 34078 15374 34130
rect 15426 34078 15428 34130
rect 15372 34066 15428 34078
rect 15484 34132 15540 36428
rect 16044 36390 16100 36428
rect 15820 36370 15876 36382
rect 15820 36318 15822 36370
rect 15874 36318 15876 36370
rect 15484 34066 15540 34076
rect 15596 36148 15652 36158
rect 15820 36148 15876 36318
rect 15652 36092 15876 36148
rect 15596 35698 15652 36092
rect 15932 35924 15988 35934
rect 16268 35924 16324 37212
rect 16380 37174 16436 37212
rect 17388 37268 17444 37326
rect 17388 37202 17444 37212
rect 16604 37154 16660 37166
rect 16604 37102 16606 37154
rect 16658 37102 16660 37154
rect 16492 37044 16548 37054
rect 16492 36372 16548 36988
rect 16604 36820 16660 37102
rect 17276 37044 17332 37054
rect 17276 36950 17332 36988
rect 16604 36764 16996 36820
rect 16940 36594 16996 36764
rect 16940 36542 16942 36594
rect 16994 36542 16996 36594
rect 16940 36530 16996 36542
rect 16716 36482 16772 36494
rect 16716 36430 16718 36482
rect 16770 36430 16772 36482
rect 16492 36316 16660 36372
rect 15932 35922 16324 35924
rect 15932 35870 15934 35922
rect 15986 35870 16324 35922
rect 15932 35868 16324 35870
rect 16380 36258 16436 36270
rect 16380 36206 16382 36258
rect 16434 36206 16436 36258
rect 15932 35858 15988 35868
rect 15708 35812 15764 35822
rect 15708 35718 15764 35756
rect 15596 35646 15598 35698
rect 15650 35646 15652 35698
rect 15148 34020 15204 34030
rect 15148 34018 15316 34020
rect 15148 33966 15150 34018
rect 15202 33966 15316 34018
rect 15148 33964 15316 33966
rect 15148 33954 15204 33964
rect 15260 33460 15316 33964
rect 15372 33460 15428 33470
rect 15316 33458 15428 33460
rect 15316 33406 15374 33458
rect 15426 33406 15428 33458
rect 15316 33404 15428 33406
rect 15260 33366 15316 33404
rect 15372 33394 15428 33404
rect 15036 33294 15038 33346
rect 15090 33294 15092 33346
rect 15036 33282 15092 33294
rect 14476 33236 14532 33246
rect 15596 33236 15652 35646
rect 16156 35476 16212 35486
rect 15708 34804 15764 34814
rect 15708 34354 15764 34748
rect 15708 34302 15710 34354
rect 15762 34302 15764 34354
rect 15708 34290 15764 34302
rect 16044 34244 16100 34254
rect 16044 34150 16100 34188
rect 16156 33572 16212 35420
rect 16380 35252 16436 36206
rect 16492 35810 16548 35822
rect 16492 35758 16494 35810
rect 16546 35758 16548 35810
rect 16492 35700 16548 35758
rect 16604 35810 16660 36316
rect 16604 35758 16606 35810
rect 16658 35758 16660 35810
rect 16604 35746 16660 35758
rect 16492 35634 16548 35644
rect 16492 35476 16548 35486
rect 16716 35476 16772 36430
rect 17164 36260 17220 36270
rect 17052 36258 17220 36260
rect 17052 36206 17166 36258
rect 17218 36206 17220 36258
rect 17052 36204 17220 36206
rect 16492 35474 16772 35476
rect 16492 35422 16494 35474
rect 16546 35422 16772 35474
rect 16492 35420 16772 35422
rect 16828 35700 16884 35710
rect 16492 35410 16548 35420
rect 16380 35196 16660 35252
rect 16268 34804 16324 34814
rect 16268 34354 16324 34748
rect 16380 34690 16436 34702
rect 16380 34638 16382 34690
rect 16434 34638 16436 34690
rect 16380 34580 16436 34638
rect 16380 34514 16436 34524
rect 16268 34302 16270 34354
rect 16322 34302 16324 34354
rect 16268 34290 16324 34302
rect 16604 34356 16660 35196
rect 16828 35028 16884 35644
rect 16828 35026 16996 35028
rect 16828 34974 16830 35026
rect 16882 34974 16996 35026
rect 16828 34972 16996 34974
rect 16828 34962 16884 34972
rect 16604 34290 16660 34300
rect 16492 34244 16548 34254
rect 16492 34150 16548 34188
rect 16604 34132 16660 34142
rect 16604 34038 16660 34076
rect 16380 34020 16436 34030
rect 16380 33926 16436 33964
rect 14252 33234 14532 33236
rect 14252 33182 14478 33234
rect 14530 33182 14532 33234
rect 14252 33180 14532 33182
rect 13580 33170 13636 33180
rect 14476 31332 14532 33180
rect 15372 33180 15652 33236
rect 15820 33458 15876 33470
rect 15820 33406 15822 33458
rect 15874 33406 15876 33458
rect 12908 31054 12910 31106
rect 12962 31054 12964 31106
rect 12908 31042 12964 31054
rect 14028 31276 14532 31332
rect 15036 31892 15204 31948
rect 12236 30942 12238 30994
rect 12290 30942 12292 30994
rect 12236 29428 12292 30942
rect 12236 29362 12292 29372
rect 12348 29986 12404 29998
rect 12348 29934 12350 29986
rect 12402 29934 12404 29986
rect 11676 29204 11732 29214
rect 11564 29148 11676 29204
rect 11676 29138 11732 29148
rect 11116 28754 11172 28812
rect 11116 28702 11118 28754
rect 11170 28702 11172 28754
rect 11116 28690 11172 28702
rect 12124 28980 12180 28990
rect 11564 28644 11620 28654
rect 11564 28550 11620 28588
rect 12012 28532 12068 28542
rect 12012 28438 12068 28476
rect 10332 27246 10334 27298
rect 10386 27246 10388 27298
rect 10332 27234 10388 27246
rect 10444 27580 10612 27636
rect 10444 26908 10500 27580
rect 10556 27412 10612 27422
rect 10556 27186 10612 27356
rect 10556 27134 10558 27186
rect 10610 27134 10612 27186
rect 10556 27122 10612 27134
rect 11004 27298 11060 27310
rect 11004 27246 11006 27298
rect 11058 27246 11060 27298
rect 11004 27186 11060 27246
rect 11004 27134 11006 27186
rect 11058 27134 11060 27186
rect 10332 26852 10500 26908
rect 11004 26908 11060 27134
rect 12124 27186 12180 28924
rect 12348 28644 12404 29934
rect 13580 29428 13636 29438
rect 13580 29334 13636 29372
rect 12908 29316 12964 29326
rect 12908 29222 12964 29260
rect 13916 29316 13972 29326
rect 13804 29092 13860 29102
rect 12348 28578 12404 28588
rect 12460 28868 12516 28878
rect 12348 28420 12404 28430
rect 12460 28420 12516 28812
rect 12572 28756 12628 28766
rect 12572 28642 12628 28700
rect 12572 28590 12574 28642
rect 12626 28590 12628 28642
rect 12572 28578 12628 28590
rect 12796 28644 12852 28654
rect 12348 28418 12516 28420
rect 12348 28366 12350 28418
rect 12402 28366 12516 28418
rect 12348 28364 12516 28366
rect 12348 28354 12404 28364
rect 12124 27134 12126 27186
rect 12178 27134 12180 27186
rect 12124 27122 12180 27134
rect 12460 27074 12516 27086
rect 12460 27022 12462 27074
rect 12514 27022 12516 27074
rect 11004 26852 11172 26908
rect 10332 25618 10388 26852
rect 10332 25566 10334 25618
rect 10386 25566 10388 25618
rect 10332 25554 10388 25566
rect 10780 25620 10836 25630
rect 10108 25506 10164 25518
rect 10108 25454 10110 25506
rect 10162 25454 10164 25506
rect 9772 24724 9828 24734
rect 10108 24724 10164 25454
rect 9772 24722 10164 24724
rect 9772 24670 9774 24722
rect 9826 24670 10164 24722
rect 9772 24668 10164 24670
rect 10220 25396 10276 25406
rect 9772 23604 9828 24668
rect 9772 23538 9828 23548
rect 9884 23380 9940 23390
rect 9884 23044 9940 23324
rect 10220 23156 10276 25340
rect 10780 24946 10836 25564
rect 10892 25396 10948 25406
rect 10892 25302 10948 25340
rect 11004 25284 11060 25294
rect 11004 25190 11060 25228
rect 11116 25060 11172 26852
rect 11452 25620 11508 25630
rect 11452 25526 11508 25564
rect 11172 25004 11284 25060
rect 11116 24994 11172 25004
rect 10780 24894 10782 24946
rect 10834 24894 10836 24946
rect 10780 24882 10836 24894
rect 10332 24836 10388 24846
rect 10332 24722 10388 24780
rect 10892 24836 10948 24846
rect 10668 24724 10724 24734
rect 10332 24670 10334 24722
rect 10386 24670 10388 24722
rect 10332 24658 10388 24670
rect 10556 24722 10724 24724
rect 10556 24670 10670 24722
rect 10722 24670 10724 24722
rect 10556 24668 10724 24670
rect 10332 23156 10388 23166
rect 10220 23154 10388 23156
rect 10220 23102 10334 23154
rect 10386 23102 10388 23154
rect 10220 23100 10388 23102
rect 10332 23090 10388 23100
rect 9772 23042 9940 23044
rect 9772 22990 9886 23042
rect 9938 22990 9940 23042
rect 9772 22988 9940 22990
rect 9548 20804 9604 20814
rect 9548 20690 9604 20748
rect 9548 20638 9550 20690
rect 9602 20638 9604 20690
rect 9548 20626 9604 20638
rect 9436 20514 9492 20524
rect 9548 20356 9604 20366
rect 9324 19684 9380 19694
rect 9212 19628 9324 19684
rect 9324 19618 9380 19628
rect 9548 19346 9604 20300
rect 9660 19908 9716 19918
rect 9772 19908 9828 22988
rect 9884 22978 9940 22988
rect 10108 20804 10164 20814
rect 10164 20748 10500 20804
rect 10108 20710 10164 20748
rect 9716 19852 9828 19908
rect 9884 20578 9940 20590
rect 9884 20526 9886 20578
rect 9938 20526 9940 20578
rect 9660 19814 9716 19852
rect 9548 19294 9550 19346
rect 9602 19294 9604 19346
rect 9548 19282 9604 19294
rect 9436 19236 9492 19246
rect 9436 18564 9492 19180
rect 9884 19236 9940 20526
rect 10332 20018 10388 20030
rect 10332 19966 10334 20018
rect 10386 19966 10388 20018
rect 9884 19170 9940 19180
rect 10108 19906 10164 19918
rect 10108 19854 10110 19906
rect 10162 19854 10164 19906
rect 9660 19124 9716 19134
rect 9660 19030 9716 19068
rect 10108 18676 10164 19854
rect 10108 18610 10164 18620
rect 9436 18498 9492 18508
rect 10332 18452 10388 19966
rect 10444 19348 10500 20748
rect 10556 20356 10612 24668
rect 10668 24658 10724 24668
rect 10780 24498 10836 24510
rect 10780 24446 10782 24498
rect 10834 24446 10836 24498
rect 10668 24052 10724 24062
rect 10780 24052 10836 24446
rect 10668 24050 10836 24052
rect 10668 23998 10670 24050
rect 10722 23998 10836 24050
rect 10668 23996 10836 23998
rect 10668 23986 10724 23996
rect 10556 20290 10612 20300
rect 10892 20132 10948 24780
rect 10892 20066 10948 20076
rect 11116 20020 11172 20030
rect 11004 19908 11060 19918
rect 10780 19906 11060 19908
rect 10780 19854 11006 19906
rect 11058 19854 11060 19906
rect 10780 19852 11060 19854
rect 10780 19458 10836 19852
rect 11004 19842 11060 19852
rect 10780 19406 10782 19458
rect 10834 19406 10836 19458
rect 10780 19394 10836 19406
rect 11116 19458 11172 19964
rect 11116 19406 11118 19458
rect 11170 19406 11172 19458
rect 11116 19394 11172 19406
rect 10556 19348 10612 19358
rect 10444 19346 10612 19348
rect 10444 19294 10558 19346
rect 10610 19294 10612 19346
rect 10444 19292 10612 19294
rect 10556 19282 10612 19292
rect 11228 19236 11284 25004
rect 11564 24724 11620 24734
rect 11452 23940 11508 23950
rect 11564 23940 11620 24668
rect 12348 24612 12404 24622
rect 12348 24518 12404 24556
rect 11452 23938 11564 23940
rect 11452 23886 11454 23938
rect 11506 23886 11564 23938
rect 11452 23884 11564 23886
rect 11452 23874 11508 23884
rect 11564 23846 11620 23884
rect 12348 23940 12404 23950
rect 12348 23154 12404 23884
rect 12348 23102 12350 23154
rect 12402 23102 12404 23154
rect 12348 23090 12404 23102
rect 11340 22484 11396 22494
rect 11340 22390 11396 22428
rect 12124 22482 12180 22494
rect 12124 22430 12126 22482
rect 12178 22430 12180 22482
rect 11676 22370 11732 22382
rect 11676 22318 11678 22370
rect 11730 22318 11732 22370
rect 11676 21812 11732 22318
rect 11676 21746 11732 21756
rect 12012 21700 12068 21710
rect 12012 21140 12068 21644
rect 11564 21084 12068 21140
rect 11340 20690 11396 20702
rect 11340 20638 11342 20690
rect 11394 20638 11396 20690
rect 11340 20468 11396 20638
rect 11564 20690 11620 21084
rect 11564 20638 11566 20690
rect 11618 20638 11620 20690
rect 11564 20626 11620 20638
rect 11676 20914 11732 20926
rect 11676 20862 11678 20914
rect 11730 20862 11732 20914
rect 11340 20402 11396 20412
rect 11676 20132 11732 20862
rect 12012 20914 12068 21084
rect 12012 20862 12014 20914
rect 12066 20862 12068 20914
rect 12012 20850 12068 20862
rect 11788 20132 11844 20142
rect 11676 20130 11844 20132
rect 11676 20078 11790 20130
rect 11842 20078 11844 20130
rect 11676 20076 11844 20078
rect 11788 20066 11844 20076
rect 12012 20132 12068 20142
rect 12124 20132 12180 22430
rect 12236 20802 12292 20814
rect 12236 20750 12238 20802
rect 12290 20750 12292 20802
rect 12236 20468 12292 20750
rect 12236 20402 12292 20412
rect 12012 20130 12180 20132
rect 12012 20078 12014 20130
rect 12066 20078 12180 20130
rect 12012 20076 12180 20078
rect 12012 20066 12068 20076
rect 12012 19906 12068 19918
rect 12012 19854 12014 19906
rect 12066 19854 12068 19906
rect 12012 19458 12068 19854
rect 12124 19908 12180 20076
rect 12236 20020 12292 20030
rect 12236 19926 12292 19964
rect 12124 19842 12180 19852
rect 12012 19406 12014 19458
rect 12066 19406 12068 19458
rect 12012 19394 12068 19406
rect 10332 18386 10388 18396
rect 10780 19180 11284 19236
rect 9100 16492 9492 16548
rect 8540 16212 8596 16222
rect 8596 16156 8708 16212
rect 8540 16118 8596 16156
rect 8316 15474 8372 15484
rect 8092 13918 8094 13970
rect 8146 13918 8148 13970
rect 7868 13858 7924 13870
rect 7868 13806 7870 13858
rect 7922 13806 7924 13858
rect 7868 12738 7924 13806
rect 8092 13412 8148 13918
rect 8204 15428 8260 15438
rect 8204 13970 8260 15372
rect 8428 15428 8484 15438
rect 8428 15334 8484 15372
rect 8540 15202 8596 15214
rect 8540 15150 8542 15202
rect 8594 15150 8596 15202
rect 8204 13918 8206 13970
rect 8258 13918 8260 13970
rect 8204 13860 8260 13918
rect 8428 14420 8484 14430
rect 8428 13970 8484 14364
rect 8540 14084 8596 15150
rect 8540 14018 8596 14028
rect 8428 13918 8430 13970
rect 8482 13918 8484 13970
rect 8428 13906 8484 13918
rect 8652 13972 8708 16156
rect 9436 16098 9492 16492
rect 9436 16046 9438 16098
rect 9490 16046 9492 16098
rect 9436 16034 9492 16046
rect 9772 15876 9828 15886
rect 9660 15874 9828 15876
rect 9660 15822 9774 15874
rect 9826 15822 9828 15874
rect 9660 15820 9828 15822
rect 9100 15540 9156 15550
rect 8988 15484 9100 15540
rect 8988 15426 9044 15484
rect 9100 15474 9156 15484
rect 8988 15374 8990 15426
rect 9042 15374 9044 15426
rect 8988 15362 9044 15374
rect 8764 15316 8820 15326
rect 9660 15316 9716 15820
rect 9772 15810 9828 15820
rect 9772 15540 9828 15578
rect 10780 15540 10836 19180
rect 12236 19122 12292 19134
rect 12236 19070 12238 19122
rect 12290 19070 12292 19122
rect 12236 18340 12292 19070
rect 12236 18274 12292 18284
rect 9772 15474 9828 15484
rect 10332 15538 10836 15540
rect 10332 15486 10782 15538
rect 10834 15486 10836 15538
rect 10332 15484 10836 15486
rect 8764 15222 8820 15260
rect 9548 15314 9716 15316
rect 9548 15262 9662 15314
rect 9714 15262 9716 15314
rect 9548 15260 9716 15262
rect 9548 15204 9604 15260
rect 9660 15250 9716 15260
rect 9772 15316 9828 15326
rect 9884 15316 9940 15326
rect 9828 15314 9940 15316
rect 9828 15262 9886 15314
rect 9938 15262 9940 15314
rect 9828 15260 9940 15262
rect 9772 15250 9828 15260
rect 8652 13906 8708 13916
rect 9100 15148 9604 15204
rect 8204 13794 8260 13804
rect 8652 13746 8708 13758
rect 8652 13694 8654 13746
rect 8706 13694 8708 13746
rect 8092 13346 8148 13356
rect 8316 13634 8372 13646
rect 8316 13582 8318 13634
rect 8370 13582 8372 13634
rect 8316 12852 8372 13582
rect 8652 13636 8708 13694
rect 9100 13636 9156 15148
rect 9436 14756 9492 14766
rect 8652 13580 9156 13636
rect 8540 13412 8596 13422
rect 8540 12964 8596 13356
rect 8652 12964 8708 12974
rect 8540 12962 8708 12964
rect 8540 12910 8654 12962
rect 8706 12910 8708 12962
rect 8540 12908 8708 12910
rect 8652 12898 8708 12908
rect 8316 12796 8596 12852
rect 7868 12686 7870 12738
rect 7922 12686 7924 12738
rect 7868 12516 7924 12686
rect 7980 12740 8036 12750
rect 7980 12646 8036 12684
rect 8092 12740 8148 12750
rect 8092 12738 8484 12740
rect 8092 12686 8094 12738
rect 8146 12686 8484 12738
rect 8092 12684 8484 12686
rect 8092 12674 8148 12684
rect 7868 12460 8036 12516
rect 7868 12180 7924 12190
rect 7812 12178 7924 12180
rect 7812 12126 7870 12178
rect 7922 12126 7924 12178
rect 7812 12124 7924 12126
rect 7756 12086 7812 12124
rect 7868 12114 7924 12124
rect 7532 11396 7588 11406
rect 7532 10834 7588 11340
rect 7980 11394 8036 12460
rect 8428 12402 8484 12684
rect 8428 12350 8430 12402
rect 8482 12350 8484 12402
rect 8428 12338 8484 12350
rect 8092 12068 8148 12078
rect 8092 11974 8148 12012
rect 8540 11620 8596 12796
rect 8764 12738 8820 12750
rect 8764 12686 8766 12738
rect 8818 12686 8820 12738
rect 8764 12404 8820 12686
rect 8764 12338 8820 12348
rect 8876 12738 8932 12750
rect 8876 12686 8878 12738
rect 8930 12686 8932 12738
rect 8540 11564 8708 11620
rect 7980 11342 7982 11394
rect 8034 11342 8036 11394
rect 7980 11330 8036 11342
rect 8428 11396 8484 11406
rect 8428 11302 8484 11340
rect 7532 10782 7534 10834
rect 7586 10782 7588 10834
rect 7532 10770 7588 10782
rect 7644 11282 7700 11294
rect 7644 11230 7646 11282
rect 7698 11230 7700 11282
rect 7644 10948 7700 11230
rect 8204 11282 8260 11294
rect 8204 11230 8206 11282
rect 8258 11230 8260 11282
rect 8204 10948 8260 11230
rect 7644 10892 8260 10948
rect 7644 10722 7700 10892
rect 8316 10836 8372 10846
rect 8316 10742 8372 10780
rect 7644 10670 7646 10722
rect 7698 10670 7700 10722
rect 7644 10658 7700 10670
rect 8204 10722 8260 10734
rect 8204 10670 8206 10722
rect 8258 10670 8260 10722
rect 7308 10558 7310 10610
rect 7362 10558 7364 10610
rect 7308 10546 7364 10558
rect 8204 10500 8260 10670
rect 8540 10722 8596 10734
rect 8540 10670 8542 10722
rect 8594 10670 8596 10722
rect 8428 10612 8484 10622
rect 8540 10612 8596 10670
rect 8428 10610 8596 10612
rect 8428 10558 8430 10610
rect 8482 10558 8596 10610
rect 8428 10556 8596 10558
rect 8428 10546 8484 10556
rect 8204 10434 8260 10444
rect 8652 10050 8708 11564
rect 8764 11396 8820 11434
rect 8764 11330 8820 11340
rect 8764 11172 8820 11182
rect 8764 11078 8820 11116
rect 8764 10836 8820 10846
rect 8876 10836 8932 12686
rect 8988 12740 9044 12750
rect 8988 12646 9044 12684
rect 9100 11284 9156 13580
rect 9212 13972 9268 13982
rect 9212 12962 9268 13916
rect 9212 12910 9214 12962
rect 9266 12910 9268 12962
rect 9212 12898 9268 12910
rect 9324 13748 9380 13758
rect 9212 11508 9268 11518
rect 9324 11508 9380 13692
rect 9212 11506 9380 11508
rect 9212 11454 9214 11506
rect 9266 11454 9380 11506
rect 9212 11452 9380 11454
rect 9436 11508 9492 14700
rect 9884 14196 9940 15260
rect 10332 15314 10388 15484
rect 10780 15474 10836 15484
rect 11564 16436 11620 16446
rect 10332 15262 10334 15314
rect 10386 15262 10388 15314
rect 10332 15250 10388 15262
rect 11564 15314 11620 16380
rect 12460 15540 12516 27022
rect 12796 26908 12852 28588
rect 13804 28642 13860 29036
rect 13804 28590 13806 28642
rect 13858 28590 13860 28642
rect 13804 28578 13860 28590
rect 13916 28642 13972 29260
rect 13916 28590 13918 28642
rect 13970 28590 13972 28642
rect 13916 28578 13972 28590
rect 13468 28532 13524 28542
rect 13468 28438 13524 28476
rect 12908 28420 12964 28430
rect 12908 27186 12964 28364
rect 13580 28420 13636 28430
rect 13580 28326 13636 28364
rect 12908 27134 12910 27186
rect 12962 27134 12964 27186
rect 12908 27122 12964 27134
rect 13356 27746 13412 27758
rect 13356 27694 13358 27746
rect 13410 27694 13412 27746
rect 12796 26852 12964 26908
rect 12572 20580 12628 20590
rect 12572 20578 12852 20580
rect 12572 20526 12574 20578
rect 12626 20526 12852 20578
rect 12572 20524 12852 20526
rect 12572 20514 12628 20524
rect 12572 20020 12628 20030
rect 12572 19926 12628 19964
rect 12796 20018 12852 20524
rect 12796 19966 12798 20018
rect 12850 19966 12852 20018
rect 12796 19954 12852 19966
rect 12908 19908 12964 26852
rect 13356 25508 13412 27694
rect 13468 25508 13524 25518
rect 13356 25506 13524 25508
rect 13356 25454 13470 25506
rect 13522 25454 13524 25506
rect 13356 25452 13524 25454
rect 13356 24724 13412 25452
rect 13468 25442 13524 25452
rect 14028 24836 14084 31276
rect 15036 30882 15092 31892
rect 15148 31826 15204 31836
rect 15036 30830 15038 30882
rect 15090 30830 15092 30882
rect 15036 30818 15092 30830
rect 14476 29316 14532 29326
rect 14140 29314 14532 29316
rect 14140 29262 14478 29314
rect 14530 29262 14532 29314
rect 14140 29260 14532 29262
rect 14140 28530 14196 29260
rect 14476 29250 14532 29260
rect 15372 28754 15428 33180
rect 15820 32564 15876 33406
rect 16044 33348 16100 33358
rect 16044 33254 16100 33292
rect 15820 31892 15876 32508
rect 15820 31798 15876 31836
rect 15932 33012 15988 33022
rect 15708 31780 15764 31790
rect 15372 28702 15374 28754
rect 15426 28702 15428 28754
rect 15372 28690 15428 28702
rect 15596 31778 15764 31780
rect 15596 31726 15710 31778
rect 15762 31726 15764 31778
rect 15596 31724 15764 31726
rect 14812 28642 14868 28654
rect 14812 28590 14814 28642
rect 14866 28590 14868 28642
rect 14140 28478 14142 28530
rect 14194 28478 14196 28530
rect 14140 28084 14196 28478
rect 14140 25620 14196 28028
rect 14252 28530 14308 28542
rect 14252 28478 14254 28530
rect 14306 28478 14308 28530
rect 14252 26964 14308 28478
rect 14812 26908 14868 28590
rect 15596 26908 15652 31724
rect 15708 31714 15764 31724
rect 15932 30994 15988 32956
rect 15932 30942 15934 30994
rect 15986 30942 15988 30994
rect 15932 30930 15988 30942
rect 16156 29652 16212 33516
rect 16828 33122 16884 33134
rect 16828 33070 16830 33122
rect 16882 33070 16884 33122
rect 16492 32564 16548 32574
rect 16828 32564 16884 33070
rect 16492 32562 16884 32564
rect 16492 32510 16494 32562
rect 16546 32510 16884 32562
rect 16492 32508 16884 32510
rect 16380 30994 16436 31006
rect 16380 30942 16382 30994
rect 16434 30942 16436 30994
rect 16380 30884 16436 30942
rect 16380 30818 16436 30828
rect 16156 29586 16212 29596
rect 15708 29428 15764 29438
rect 15708 28644 15764 29372
rect 16156 29204 16212 29214
rect 16156 28644 16212 29148
rect 15708 28642 15876 28644
rect 15708 28590 15710 28642
rect 15762 28590 15876 28642
rect 15708 28588 15876 28590
rect 15708 28578 15764 28588
rect 15820 27188 15876 28588
rect 15932 27860 15988 27870
rect 15932 27766 15988 27804
rect 15932 27188 15988 27198
rect 15820 27186 15988 27188
rect 15820 27134 15934 27186
rect 15986 27134 15988 27186
rect 15820 27132 15988 27134
rect 15932 27122 15988 27132
rect 16156 27074 16212 28588
rect 16380 27860 16436 27870
rect 16492 27860 16548 32508
rect 16940 31892 16996 34972
rect 16940 31826 16996 31836
rect 17052 33236 17108 36204
rect 17164 36194 17220 36204
rect 17276 36258 17332 36270
rect 17276 36206 17278 36258
rect 17330 36206 17332 36258
rect 17276 35812 17332 36206
rect 17388 36260 17444 36270
rect 17388 36258 17668 36260
rect 17388 36206 17390 36258
rect 17442 36206 17668 36258
rect 17388 36204 17668 36206
rect 17388 36194 17444 36204
rect 17388 35812 17444 35822
rect 17276 35810 17444 35812
rect 17276 35758 17390 35810
rect 17442 35758 17444 35810
rect 17276 35756 17444 35758
rect 17388 35746 17444 35756
rect 17500 35810 17556 35822
rect 17500 35758 17502 35810
rect 17554 35758 17556 35810
rect 17500 35364 17556 35758
rect 17500 35298 17556 35308
rect 17612 34580 17668 36204
rect 17724 35922 17780 37884
rect 18396 37874 18452 37884
rect 19180 37828 19236 37998
rect 21420 37940 21476 37950
rect 21420 37846 21476 37884
rect 21644 37938 21700 37950
rect 21644 37886 21646 37938
rect 21698 37886 21700 37938
rect 19628 37828 19684 37838
rect 19180 37826 19684 37828
rect 19180 37774 19630 37826
rect 19682 37774 19684 37826
rect 19180 37772 19684 37774
rect 19628 37492 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37436 19908 37492
rect 17836 37266 17892 37278
rect 17836 37214 17838 37266
rect 17890 37214 17892 37266
rect 17836 37156 17892 37214
rect 17836 37090 17892 37100
rect 19628 37154 19684 37166
rect 19628 37102 19630 37154
rect 19682 37102 19684 37154
rect 17836 36484 17892 36494
rect 17836 36390 17892 36428
rect 19404 36484 19460 36494
rect 19628 36484 19684 37102
rect 19852 37044 19908 37436
rect 19852 36978 19908 36988
rect 19404 36482 19684 36484
rect 19404 36430 19406 36482
rect 19458 36430 19684 36482
rect 19404 36428 19684 36430
rect 20188 36482 20244 36494
rect 20188 36430 20190 36482
rect 20242 36430 20244 36482
rect 18956 36370 19012 36382
rect 18956 36318 18958 36370
rect 19010 36318 19012 36370
rect 17724 35870 17726 35922
rect 17778 35870 17780 35922
rect 17724 35858 17780 35870
rect 18172 36258 18228 36270
rect 18172 36206 18174 36258
rect 18226 36206 18228 36258
rect 18060 35586 18116 35598
rect 18060 35534 18062 35586
rect 18114 35534 18116 35586
rect 18060 35364 18116 35534
rect 18060 35298 18116 35308
rect 17612 34514 17668 34524
rect 16604 31780 16660 31790
rect 16604 31686 16660 31724
rect 16828 30884 16884 30894
rect 16716 30882 16884 30884
rect 16716 30830 16830 30882
rect 16882 30830 16884 30882
rect 16716 30828 16884 30830
rect 16716 30212 16772 30828
rect 16828 30818 16884 30828
rect 16716 30146 16772 30156
rect 16716 29876 16772 29886
rect 16604 29820 16716 29876
rect 16604 29204 16660 29820
rect 16716 29810 16772 29820
rect 16716 29652 16772 29662
rect 16716 29558 16772 29596
rect 16940 29540 16996 29550
rect 16828 29428 16884 29438
rect 16940 29428 16996 29484
rect 16828 29426 16996 29428
rect 16828 29374 16830 29426
rect 16882 29374 16996 29426
rect 16828 29372 16996 29374
rect 16828 29362 16884 29372
rect 16716 29204 16772 29214
rect 16604 29202 16772 29204
rect 16604 29150 16718 29202
rect 16770 29150 16772 29202
rect 16604 29148 16772 29150
rect 16716 29138 16772 29148
rect 17052 28754 17108 33180
rect 17052 28702 17054 28754
rect 17106 28702 17108 28754
rect 17052 28690 17108 28702
rect 17164 33348 17220 33358
rect 18172 33348 18228 36206
rect 18956 35812 19012 36318
rect 18844 34802 18900 34814
rect 18844 34750 18846 34802
rect 18898 34750 18900 34802
rect 18844 34132 18900 34750
rect 18956 34802 19012 35756
rect 19404 35700 19460 36428
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19404 35634 19460 35644
rect 20188 35588 20244 36430
rect 20748 36484 20804 36494
rect 20972 36484 21028 36494
rect 21532 36484 21588 36494
rect 20748 36482 20972 36484
rect 20748 36430 20750 36482
rect 20802 36430 20972 36482
rect 20748 36428 20972 36430
rect 20748 36418 20804 36428
rect 20972 36418 21028 36428
rect 21084 36482 21588 36484
rect 21084 36430 21534 36482
rect 21586 36430 21588 36482
rect 21084 36428 21588 36430
rect 20860 35924 20916 35934
rect 21084 35924 21140 36428
rect 21532 36418 21588 36428
rect 21644 36482 21700 37886
rect 21756 37378 21812 38108
rect 23212 37940 23268 38780
rect 23212 37490 23268 37884
rect 23212 37438 23214 37490
rect 23266 37438 23268 37490
rect 23212 37426 23268 37438
rect 21756 37326 21758 37378
rect 21810 37326 21812 37378
rect 21756 37314 21812 37326
rect 22540 37266 22596 37278
rect 22540 37214 22542 37266
rect 22594 37214 22596 37266
rect 22540 37044 22596 37214
rect 22540 36978 22596 36988
rect 22876 37266 22932 37278
rect 22876 37214 22878 37266
rect 22930 37214 22932 37266
rect 21644 36430 21646 36482
rect 21698 36430 21700 36482
rect 21644 36418 21700 36430
rect 21756 36484 21812 36494
rect 21756 36390 21812 36428
rect 21868 36482 21924 36494
rect 21868 36430 21870 36482
rect 21922 36430 21924 36482
rect 21868 36372 21924 36430
rect 21868 36306 21924 36316
rect 21420 36260 21476 36270
rect 22540 36260 22596 36270
rect 22876 36260 22932 37214
rect 23436 37044 23492 37054
rect 23548 37044 23604 39340
rect 25340 39058 25396 39452
rect 25340 39006 25342 39058
rect 25394 39006 25396 39058
rect 25340 38994 25396 39006
rect 25564 39508 25620 39518
rect 25564 38836 25620 39452
rect 25564 38742 25620 38780
rect 25228 38724 25284 38734
rect 25116 38722 25284 38724
rect 25116 38670 25230 38722
rect 25282 38670 25284 38722
rect 25116 38668 25284 38670
rect 25116 38162 25172 38668
rect 25228 38658 25284 38668
rect 26124 38668 26180 39676
rect 26348 39666 26404 39676
rect 26796 39396 26852 40348
rect 29148 40404 29204 40414
rect 29372 40404 29428 40910
rect 30268 40962 30436 40964
rect 30268 40910 30382 40962
rect 30434 40910 30436 40962
rect 30268 40908 30436 40910
rect 29596 40404 29652 40414
rect 29372 40348 29596 40404
rect 29148 40310 29204 40348
rect 29596 40310 29652 40348
rect 27244 40292 27300 40302
rect 27244 39842 27300 40236
rect 27244 39790 27246 39842
rect 27298 39790 27300 39842
rect 27244 39778 27300 39790
rect 28700 40290 28756 40302
rect 28700 40238 28702 40290
rect 28754 40238 28756 40290
rect 28700 39620 28756 40238
rect 29372 39620 29428 39630
rect 28700 39618 29428 39620
rect 28700 39566 29374 39618
rect 29426 39566 29428 39618
rect 28700 39564 29428 39566
rect 27356 39508 27412 39518
rect 27356 39414 27412 39452
rect 27580 39508 27636 39518
rect 27580 39506 28084 39508
rect 27580 39454 27582 39506
rect 27634 39454 28084 39506
rect 27580 39452 28084 39454
rect 27580 39442 27636 39452
rect 26796 39302 26852 39340
rect 27916 38724 27972 38734
rect 26124 38612 26628 38668
rect 25116 38110 25118 38162
rect 25170 38110 25172 38162
rect 25116 38098 25172 38110
rect 26572 38164 26628 38612
rect 27468 38612 27972 38668
rect 26572 38108 26852 38164
rect 25340 38050 25396 38062
rect 25340 37998 25342 38050
rect 25394 37998 25396 38050
rect 24668 37938 24724 37950
rect 24668 37886 24670 37938
rect 24722 37886 24724 37938
rect 23660 37154 23716 37166
rect 23660 37102 23662 37154
rect 23714 37102 23716 37154
rect 23660 37044 23716 37102
rect 23492 36988 23716 37044
rect 21420 36258 21700 36260
rect 21420 36206 21422 36258
rect 21474 36206 21700 36258
rect 21420 36204 21700 36206
rect 21420 36194 21476 36204
rect 19740 35532 20244 35588
rect 20300 35922 21140 35924
rect 20300 35870 20862 35922
rect 20914 35870 21140 35922
rect 20300 35868 21140 35870
rect 19740 34914 19796 35532
rect 19740 34862 19742 34914
rect 19794 34862 19796 34914
rect 19740 34850 19796 34862
rect 18956 34750 18958 34802
rect 19010 34750 19012 34802
rect 18956 34738 19012 34750
rect 19404 34804 19460 34814
rect 19404 34710 19460 34748
rect 19180 34692 19236 34702
rect 19180 34690 19348 34692
rect 19180 34638 19182 34690
rect 19234 34638 19348 34690
rect 19180 34636 19348 34638
rect 19180 34626 19236 34636
rect 19292 34580 19348 34636
rect 19516 34690 19572 34702
rect 19516 34638 19518 34690
rect 19570 34638 19572 34690
rect 19516 34580 19572 34638
rect 19292 34524 19572 34580
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 20188 34356 20244 34366
rect 19516 34244 19572 34254
rect 19516 34150 19572 34188
rect 19852 34244 19908 34254
rect 19180 34132 19236 34142
rect 19740 34132 19796 34142
rect 18844 34130 19236 34132
rect 18844 34078 19182 34130
rect 19234 34078 19236 34130
rect 18844 34076 19236 34078
rect 18620 33572 18676 33582
rect 18620 33478 18676 33516
rect 18396 33348 18452 33358
rect 18172 33346 18452 33348
rect 18172 33294 18398 33346
rect 18450 33294 18452 33346
rect 18172 33292 18452 33294
rect 17164 32004 17220 33292
rect 18396 33236 18452 33292
rect 18396 33170 18452 33180
rect 18956 33122 19012 33134
rect 18956 33070 18958 33122
rect 19010 33070 19012 33122
rect 18956 32788 19012 33070
rect 18732 32732 18956 32788
rect 17724 32674 17780 32686
rect 17724 32622 17726 32674
rect 17778 32622 17780 32674
rect 17388 32564 17444 32574
rect 17388 32470 17444 32508
rect 17724 32340 17780 32622
rect 17724 32274 17780 32284
rect 18396 32564 18452 32574
rect 16436 27804 16548 27860
rect 16828 28642 16884 28654
rect 16828 28590 16830 28642
rect 16882 28590 16884 28642
rect 16380 27766 16436 27804
rect 16828 27636 16884 28590
rect 16156 27022 16158 27074
rect 16210 27022 16212 27074
rect 16156 27010 16212 27022
rect 16380 27580 16884 27636
rect 14252 26898 14308 26908
rect 14140 25554 14196 25564
rect 14476 26852 14868 26908
rect 15484 26852 15652 26908
rect 14028 24770 14084 24780
rect 14252 25394 14308 25406
rect 14252 25342 14254 25394
rect 14306 25342 14308 25394
rect 13356 24658 13412 24668
rect 14252 23828 14308 25342
rect 14252 23762 14308 23772
rect 14476 24610 14532 26852
rect 14476 24558 14478 24610
rect 14530 24558 14532 24610
rect 13020 23156 13076 23166
rect 13020 23062 13076 23100
rect 14476 21924 14532 24558
rect 15484 23268 15540 26852
rect 16380 25620 16436 27580
rect 17164 27298 17220 31948
rect 18172 31780 18228 31790
rect 17500 30884 17556 30894
rect 17500 29764 17556 30828
rect 17164 27246 17166 27298
rect 17218 27246 17220 27298
rect 17164 27234 17220 27246
rect 17276 29708 17556 29764
rect 17836 30210 17892 30222
rect 17836 30158 17838 30210
rect 17890 30158 17892 30210
rect 16716 27188 16772 27198
rect 16716 27076 16772 27132
rect 16828 27076 16884 27086
rect 16716 27074 16884 27076
rect 16716 27022 16830 27074
rect 16882 27022 16884 27074
rect 16716 27020 16884 27022
rect 16828 27010 16884 27020
rect 17276 26908 17332 29708
rect 17500 29540 17556 29550
rect 17556 29484 17668 29540
rect 17500 29446 17556 29484
rect 17388 29428 17444 29438
rect 17388 29334 17444 29372
rect 17500 29204 17556 29214
rect 17500 29110 17556 29148
rect 17500 28868 17556 28878
rect 17388 28812 17500 28868
rect 17388 28084 17444 28812
rect 17500 28802 17556 28812
rect 17612 28532 17668 29484
rect 17836 28868 17892 30158
rect 17948 30212 18004 30222
rect 17948 30118 18004 30156
rect 18172 30210 18228 31724
rect 18172 30158 18174 30210
rect 18226 30158 18228 30210
rect 18172 30146 18228 30158
rect 18284 30772 18340 30782
rect 18284 29426 18340 30716
rect 18396 30210 18452 32508
rect 18620 32564 18676 32574
rect 18732 32564 18788 32732
rect 18956 32694 19012 32732
rect 19068 32674 19124 34076
rect 19180 34066 19236 34076
rect 19628 34076 19740 34132
rect 19292 33572 19348 33582
rect 19292 33346 19348 33516
rect 19292 33294 19294 33346
rect 19346 33294 19348 33346
rect 19292 33282 19348 33294
rect 19628 33290 19684 34076
rect 19740 34066 19796 34076
rect 19516 33236 19572 33246
rect 19628 33238 19630 33290
rect 19682 33238 19684 33290
rect 19628 33226 19684 33238
rect 19852 33236 19908 34188
rect 20188 34130 20244 34300
rect 20188 34078 20190 34130
rect 20242 34078 20244 34130
rect 20188 34066 20244 34078
rect 20300 34132 20356 35868
rect 20860 35858 20916 35868
rect 19740 33234 19908 33236
rect 19516 33142 19572 33180
rect 19740 33182 19854 33234
rect 19906 33182 19908 33234
rect 19740 33180 19908 33182
rect 19740 33124 19796 33180
rect 19852 33170 19908 33180
rect 20076 33458 20132 33470
rect 20076 33406 20078 33458
rect 20130 33406 20132 33458
rect 19068 32622 19070 32674
rect 19122 32622 19124 32674
rect 18620 32562 18788 32564
rect 18620 32510 18622 32562
rect 18674 32510 18788 32562
rect 18620 32508 18788 32510
rect 18844 32564 18900 32574
rect 18620 31892 18676 32508
rect 18844 32470 18900 32508
rect 19068 32340 19124 32622
rect 19628 33068 19796 33124
rect 20076 33124 20132 33406
rect 20076 33068 20244 33124
rect 19628 32674 19684 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32622 19630 32674
rect 19682 32622 19684 32674
rect 19628 32610 19684 32622
rect 19740 32788 19796 32798
rect 20188 32788 20244 33068
rect 19796 32732 20020 32788
rect 19404 32564 19460 32574
rect 19404 32470 19460 32508
rect 19068 32274 19124 32284
rect 19180 32340 19236 32350
rect 19180 32338 19348 32340
rect 19180 32286 19182 32338
rect 19234 32286 19348 32338
rect 19180 32284 19348 32286
rect 19180 32274 19236 32284
rect 18732 31892 18788 31902
rect 18620 31890 18788 31892
rect 18620 31838 18734 31890
rect 18786 31838 18788 31890
rect 18620 31836 18788 31838
rect 18732 31826 18788 31836
rect 18508 31780 18564 31790
rect 18508 31686 18564 31724
rect 19180 31666 19236 31678
rect 19180 31614 19182 31666
rect 19234 31614 19236 31666
rect 19068 31220 19124 31230
rect 19180 31220 19236 31614
rect 19068 31218 19236 31220
rect 19068 31166 19070 31218
rect 19122 31166 19236 31218
rect 19068 31164 19236 31166
rect 19068 31154 19124 31164
rect 19180 30996 19236 31006
rect 19292 30996 19348 32284
rect 19740 31778 19796 32732
rect 19964 32562 20020 32732
rect 19964 32510 19966 32562
rect 20018 32510 20020 32562
rect 19964 32498 20020 32510
rect 20076 32732 20244 32788
rect 19852 32450 19908 32462
rect 19852 32398 19854 32450
rect 19906 32398 19908 32450
rect 19852 31892 19908 32398
rect 19852 31826 19908 31836
rect 19740 31726 19742 31778
rect 19794 31726 19796 31778
rect 19740 31714 19796 31726
rect 20076 31780 20132 32732
rect 20300 32564 20356 34076
rect 20076 31714 20132 31724
rect 20188 32508 20356 32564
rect 20412 35700 20468 35710
rect 20524 35700 20580 35710
rect 20468 35698 20580 35700
rect 20468 35646 20526 35698
rect 20578 35646 20580 35698
rect 20468 35644 20580 35646
rect 20412 32564 20468 35644
rect 20524 35634 20580 35644
rect 20524 34244 20580 34254
rect 20524 34130 20580 34188
rect 20524 34078 20526 34130
rect 20578 34078 20580 34130
rect 20524 34066 20580 34078
rect 21532 34020 21588 34030
rect 21644 34020 21700 36204
rect 22540 36258 22932 36260
rect 22540 36206 22542 36258
rect 22594 36206 22932 36258
rect 22540 36204 22932 36206
rect 23324 36372 23380 36382
rect 21588 33964 22148 34020
rect 21532 33954 21588 33964
rect 20636 33906 20692 33918
rect 20636 33854 20638 33906
rect 20690 33854 20692 33906
rect 20636 32788 20692 33854
rect 22092 33234 22148 33964
rect 22092 33182 22094 33234
rect 22146 33182 22148 33234
rect 22092 33170 22148 33182
rect 20636 32722 20692 32732
rect 22428 33122 22484 33134
rect 22428 33070 22430 33122
rect 22482 33070 22484 33122
rect 20524 32564 20580 32574
rect 20412 32562 20580 32564
rect 20412 32510 20526 32562
rect 20578 32510 20580 32562
rect 20412 32508 20580 32510
rect 20076 31556 20132 31566
rect 20188 31556 20244 32508
rect 20524 32498 20580 32508
rect 20636 32564 20692 32574
rect 20300 32340 20356 32350
rect 20300 31666 20356 32284
rect 20636 32338 20692 32508
rect 20636 32286 20638 32338
rect 20690 32286 20692 32338
rect 20636 32274 20692 32286
rect 20748 32562 20804 32574
rect 20748 32510 20750 32562
rect 20802 32510 20804 32562
rect 20748 32116 20804 32510
rect 20300 31614 20302 31666
rect 20354 31614 20356 31666
rect 20300 31602 20356 31614
rect 20524 32060 20804 32116
rect 20076 31554 20244 31556
rect 20076 31502 20078 31554
rect 20130 31502 20244 31554
rect 20076 31500 20244 31502
rect 20412 31554 20468 31566
rect 20412 31502 20414 31554
rect 20466 31502 20468 31554
rect 20076 31490 20132 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19180 30994 19348 30996
rect 19180 30942 19182 30994
rect 19234 30942 19348 30994
rect 19180 30940 19348 30942
rect 19180 30930 19236 30940
rect 19068 30772 19124 30782
rect 19068 30678 19124 30716
rect 18396 30158 18398 30210
rect 18450 30158 18452 30210
rect 18396 30146 18452 30158
rect 18732 30212 18788 30222
rect 18732 30098 18788 30156
rect 18732 30046 18734 30098
rect 18786 30046 18788 30098
rect 18732 30034 18788 30046
rect 19180 30098 19236 30110
rect 19180 30046 19182 30098
rect 19234 30046 19236 30098
rect 18508 29988 18564 29998
rect 18508 29894 18564 29932
rect 18620 29986 18676 29998
rect 18956 29988 19012 29998
rect 18620 29934 18622 29986
rect 18674 29934 18676 29986
rect 18284 29374 18286 29426
rect 18338 29374 18340 29426
rect 18284 29362 18340 29374
rect 18396 29652 18452 29662
rect 18060 29314 18116 29326
rect 18060 29262 18062 29314
rect 18114 29262 18116 29314
rect 18060 29092 18116 29262
rect 18060 29026 18116 29036
rect 17836 28812 18116 28868
rect 17724 28532 17780 28542
rect 17612 28530 17780 28532
rect 17612 28478 17726 28530
rect 17778 28478 17780 28530
rect 17612 28476 17780 28478
rect 17388 28028 17668 28084
rect 17500 27860 17556 27870
rect 16940 26852 17332 26908
rect 17388 27858 17556 27860
rect 17388 27806 17502 27858
rect 17554 27806 17556 27858
rect 17388 27804 17556 27806
rect 17388 26852 17444 27804
rect 17500 27794 17556 27804
rect 17612 27746 17668 28028
rect 17612 27694 17614 27746
rect 17666 27694 17668 27746
rect 17612 27682 17668 27694
rect 17724 27748 17780 28476
rect 17836 27970 17892 28812
rect 18060 28754 18116 28812
rect 18060 28702 18062 28754
rect 18114 28702 18116 28754
rect 18060 28690 18116 28702
rect 18172 28644 18228 28654
rect 18172 28550 18228 28588
rect 18396 28082 18452 29596
rect 18508 29428 18564 29438
rect 18620 29428 18676 29934
rect 18508 29426 18676 29428
rect 18508 29374 18510 29426
rect 18562 29374 18676 29426
rect 18508 29372 18676 29374
rect 18844 29986 19012 29988
rect 18844 29934 18958 29986
rect 19010 29934 19012 29986
rect 18844 29932 19012 29934
rect 18508 29362 18564 29372
rect 18844 28868 18900 29932
rect 18956 29922 19012 29932
rect 19180 29876 19236 30046
rect 19180 29810 19236 29820
rect 19404 29988 19460 29998
rect 18956 29652 19012 29662
rect 18956 29650 19348 29652
rect 18956 29598 18958 29650
rect 19010 29598 19348 29650
rect 18956 29596 19348 29598
rect 18956 29586 19012 29596
rect 19292 29538 19348 29596
rect 19292 29486 19294 29538
rect 19346 29486 19348 29538
rect 19292 29474 19348 29486
rect 19180 29428 19236 29438
rect 18844 28802 18900 28812
rect 18956 29426 19236 29428
rect 18956 29374 19182 29426
rect 19234 29374 19236 29426
rect 18956 29372 19236 29374
rect 18396 28030 18398 28082
rect 18450 28030 18452 28082
rect 18396 28018 18452 28030
rect 18732 28642 18788 28654
rect 18732 28590 18734 28642
rect 18786 28590 18788 28642
rect 17836 27918 17838 27970
rect 17890 27918 17892 27970
rect 17836 27906 17892 27918
rect 18508 27970 18564 27982
rect 18508 27918 18510 27970
rect 18562 27918 18564 27970
rect 18172 27860 18228 27870
rect 17948 27858 18228 27860
rect 17948 27806 18174 27858
rect 18226 27806 18228 27858
rect 17948 27804 18228 27806
rect 17948 27748 18004 27804
rect 18172 27794 18228 27804
rect 17724 27692 18004 27748
rect 18284 27186 18340 27198
rect 18284 27134 18286 27186
rect 18338 27134 18340 27186
rect 17500 27076 17556 27086
rect 18284 27076 18340 27134
rect 18508 27188 18564 27918
rect 18732 27748 18788 28590
rect 18732 27682 18788 27692
rect 18844 27858 18900 27870
rect 18844 27806 18846 27858
rect 18898 27806 18900 27858
rect 18508 27122 18564 27132
rect 17500 27074 18340 27076
rect 17500 27022 17502 27074
rect 17554 27022 18340 27074
rect 17500 27020 18340 27022
rect 17500 27010 17556 27020
rect 18396 26962 18452 26974
rect 18396 26910 18398 26962
rect 18450 26910 18452 26962
rect 17612 26852 17668 26862
rect 16380 25618 16660 25620
rect 16380 25566 16382 25618
rect 16434 25566 16660 25618
rect 16380 25564 16660 25566
rect 16380 25554 16436 25564
rect 16604 23940 16660 25564
rect 16492 23938 16660 23940
rect 16492 23886 16606 23938
rect 16658 23886 16660 23938
rect 16492 23884 16660 23886
rect 16380 23716 16436 23726
rect 16380 23622 16436 23660
rect 15484 23174 15540 23212
rect 16380 23268 16436 23278
rect 16380 23174 16436 23212
rect 15820 23154 15876 23166
rect 15820 23102 15822 23154
rect 15874 23102 15876 23154
rect 15148 23042 15204 23054
rect 15148 22990 15150 23042
rect 15202 22990 15204 23042
rect 15148 22932 15204 22990
rect 15820 22932 15876 23102
rect 16268 23156 16324 23166
rect 16268 23062 16324 23100
rect 16156 23044 16212 23054
rect 15148 22876 15876 22932
rect 15708 22596 15764 22606
rect 15708 22482 15764 22540
rect 15708 22430 15710 22482
rect 15762 22430 15764 22482
rect 14476 21858 14532 21868
rect 15372 22370 15428 22382
rect 15372 22318 15374 22370
rect 15426 22318 15428 22370
rect 13916 21700 13972 21710
rect 13916 21606 13972 21644
rect 15372 21700 15428 22318
rect 15372 21606 15428 21644
rect 15708 21698 15764 22430
rect 15820 22148 15876 22876
rect 15932 23042 16212 23044
rect 15932 22990 16158 23042
rect 16210 22990 16212 23042
rect 15932 22988 16212 22990
rect 15932 22370 15988 22988
rect 16156 22978 16212 22988
rect 16492 22594 16548 23884
rect 16604 23874 16660 23884
rect 16828 23940 16884 23950
rect 16828 23716 16884 23884
rect 16716 22596 16772 22606
rect 16492 22542 16494 22594
rect 16546 22542 16548 22594
rect 16268 22372 16324 22382
rect 15932 22318 15934 22370
rect 15986 22318 15988 22370
rect 15932 22306 15988 22318
rect 16044 22370 16324 22372
rect 16044 22318 16270 22370
rect 16322 22318 16324 22370
rect 16044 22316 16324 22318
rect 16044 22148 16100 22316
rect 16268 22306 16324 22316
rect 15820 22092 16100 22148
rect 15708 21646 15710 21698
rect 15762 21646 15764 21698
rect 15708 21634 15764 21646
rect 16044 21924 16100 21934
rect 13580 21586 13636 21598
rect 13580 21534 13582 21586
rect 13634 21534 13636 21586
rect 13580 21364 13636 21534
rect 15260 21588 15316 21598
rect 15260 21494 15316 21532
rect 15596 21476 15652 21486
rect 15596 21382 15652 21420
rect 13468 20690 13524 20702
rect 13468 20638 13470 20690
rect 13522 20638 13524 20690
rect 13468 20468 13524 20638
rect 13580 20690 13636 21308
rect 13580 20638 13582 20690
rect 13634 20638 13636 20690
rect 13580 20626 13636 20638
rect 16044 20690 16100 21868
rect 16380 21700 16436 21710
rect 16492 21700 16548 22542
rect 16380 21698 16548 21700
rect 16380 21646 16382 21698
rect 16434 21646 16548 21698
rect 16380 21644 16548 21646
rect 16604 22540 16716 22596
rect 16380 21634 16436 21644
rect 16156 21588 16212 21598
rect 16156 21494 16212 21532
rect 16268 21586 16324 21598
rect 16268 21534 16270 21586
rect 16322 21534 16324 21586
rect 16268 21364 16324 21534
rect 16268 21298 16324 21308
rect 16604 21028 16660 22540
rect 16716 22530 16772 22540
rect 16716 22370 16772 22382
rect 16716 22318 16718 22370
rect 16770 22318 16772 22370
rect 16716 21924 16772 22318
rect 16716 21858 16772 21868
rect 16828 21700 16884 23660
rect 16716 21644 16884 21700
rect 16716 21252 16772 21644
rect 16940 21588 16996 26852
rect 17388 26850 17668 26852
rect 17388 26798 17614 26850
rect 17666 26798 17668 26850
rect 17388 26796 17668 26798
rect 17612 26516 17668 26796
rect 17724 26852 17780 26862
rect 17724 26758 17780 26796
rect 17836 26852 18340 26908
rect 17836 26850 17892 26852
rect 17836 26798 17838 26850
rect 17890 26798 17892 26850
rect 17836 26786 17892 26798
rect 17612 26450 17668 26460
rect 18284 26292 18340 26852
rect 18396 26516 18452 26910
rect 18396 26450 18452 26460
rect 18620 26962 18676 26974
rect 18620 26910 18622 26962
rect 18674 26910 18676 26962
rect 18620 26404 18676 26910
rect 18844 26740 18900 27806
rect 18956 27746 19012 29372
rect 19180 29362 19236 29372
rect 19404 28642 19460 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20412 29428 20468 31502
rect 20412 29362 20468 29372
rect 20076 29314 20132 29326
rect 20076 29262 20078 29314
rect 20130 29262 20132 29314
rect 19852 29204 19908 29214
rect 19628 29092 19684 29102
rect 19628 28866 19684 29036
rect 19628 28814 19630 28866
rect 19682 28814 19684 28866
rect 19628 28802 19684 28814
rect 19852 28866 19908 29148
rect 19852 28814 19854 28866
rect 19906 28814 19908 28866
rect 19852 28802 19908 28814
rect 19404 28590 19406 28642
rect 19458 28590 19460 28642
rect 19404 28578 19460 28590
rect 19516 28420 19572 28430
rect 20076 28420 20132 29262
rect 19516 28418 19684 28420
rect 19516 28366 19518 28418
rect 19570 28366 19684 28418
rect 19516 28364 19684 28366
rect 20076 28364 20244 28420
rect 19516 28354 19572 28364
rect 18956 27694 18958 27746
rect 19010 27694 19012 27746
rect 18956 27682 19012 27694
rect 19404 27748 19460 27758
rect 18732 26684 18900 26740
rect 19292 27188 19348 27198
rect 19292 27074 19348 27132
rect 19292 27022 19294 27074
rect 19346 27022 19348 27074
rect 18732 26516 18788 26684
rect 19180 26516 19236 26526
rect 18732 26460 18900 26516
rect 18620 26348 18788 26404
rect 18284 26236 18676 26292
rect 18508 25060 18564 25070
rect 17500 24722 17556 24734
rect 17500 24670 17502 24722
rect 17554 24670 17556 24722
rect 17052 23940 17108 23950
rect 17052 23846 17108 23884
rect 17276 23940 17332 23950
rect 17500 23940 17556 24670
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17612 24612 17668 24622
rect 17612 24518 17668 24556
rect 17836 24164 17892 24670
rect 17836 24098 17892 24108
rect 18060 24722 18116 24734
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 18060 24050 18116 24670
rect 18060 23998 18062 24050
rect 18114 23998 18116 24050
rect 18060 23986 18116 23998
rect 18508 24052 18564 25004
rect 17724 23940 17780 23950
rect 18172 23940 18228 23950
rect 17500 23938 17892 23940
rect 17500 23886 17726 23938
rect 17778 23886 17892 23938
rect 17500 23884 17892 23886
rect 17276 23846 17332 23884
rect 17724 23874 17780 23884
rect 17500 23714 17556 23726
rect 17500 23662 17502 23714
rect 17554 23662 17556 23714
rect 17500 23268 17556 23662
rect 17836 23716 17892 23884
rect 18060 23828 18116 23838
rect 17948 23716 18004 23726
rect 17836 23714 18004 23716
rect 17836 23662 17950 23714
rect 18002 23662 18004 23714
rect 17836 23660 18004 23662
rect 17500 23212 17780 23268
rect 17724 23154 17780 23212
rect 17724 23102 17726 23154
rect 17778 23102 17780 23154
rect 17724 23090 17780 23102
rect 17612 22930 17668 22942
rect 17612 22878 17614 22930
rect 17666 22878 17668 22930
rect 17612 22596 17668 22878
rect 17612 22530 17668 22540
rect 17836 22260 17892 23660
rect 17948 23650 18004 23660
rect 18060 23266 18116 23772
rect 18172 23716 18228 23884
rect 18508 23938 18564 23996
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18508 23874 18564 23886
rect 18228 23660 18340 23716
rect 18172 23622 18228 23660
rect 18060 23214 18062 23266
rect 18114 23214 18116 23266
rect 18060 23202 18116 23214
rect 17948 23156 18004 23166
rect 17948 23062 18004 23100
rect 17612 22204 17892 22260
rect 18284 22258 18340 23660
rect 18508 23156 18564 23166
rect 18508 23062 18564 23100
rect 18284 22206 18286 22258
rect 18338 22206 18340 22258
rect 17164 22146 17220 22158
rect 17164 22094 17166 22146
rect 17218 22094 17220 22146
rect 17164 21812 17220 22094
rect 17500 21812 17556 21822
rect 17164 21756 17500 21812
rect 17500 21746 17556 21756
rect 16940 21532 17220 21588
rect 16828 21474 16884 21486
rect 16828 21422 16830 21474
rect 16882 21422 16884 21474
rect 16828 21364 16884 21422
rect 17052 21364 17108 21374
rect 16828 21308 17052 21364
rect 17052 21298 17108 21308
rect 16716 21196 16884 21252
rect 16828 21140 16884 21196
rect 16828 21074 16884 21084
rect 16716 21028 16772 21038
rect 16604 21026 16772 21028
rect 16604 20974 16718 21026
rect 16770 20974 16772 21026
rect 16604 20972 16772 20974
rect 16716 20962 16772 20972
rect 17164 20916 17220 21532
rect 16940 20860 17220 20916
rect 17388 21140 17444 21150
rect 16044 20638 16046 20690
rect 16098 20638 16100 20690
rect 13468 20402 13524 20412
rect 13804 20578 13860 20590
rect 13804 20526 13806 20578
rect 13858 20526 13860 20578
rect 13804 20244 13860 20526
rect 13804 20178 13860 20188
rect 13132 20132 13188 20142
rect 13132 20038 13188 20076
rect 13356 20130 13412 20142
rect 13356 20078 13358 20130
rect 13410 20078 13412 20130
rect 13356 19908 13412 20078
rect 13916 20130 13972 20142
rect 13916 20078 13918 20130
rect 13970 20078 13972 20130
rect 12908 19852 13188 19908
rect 12796 19460 12852 19470
rect 12796 19366 12852 19404
rect 12572 19236 12628 19246
rect 12572 19142 12628 19180
rect 12908 19012 12964 19022
rect 12908 19010 13076 19012
rect 12908 18958 12910 19010
rect 12962 18958 13076 19010
rect 12908 18956 13076 18958
rect 12908 18946 12964 18956
rect 12908 18562 12964 18574
rect 12908 18510 12910 18562
rect 12962 18510 12964 18562
rect 12796 18452 12852 18462
rect 12908 18452 12964 18510
rect 12852 18396 12964 18452
rect 12796 18386 12852 18396
rect 12908 18116 12964 18396
rect 13020 18452 13076 18956
rect 13020 18386 13076 18396
rect 12908 18050 12964 18060
rect 12460 15474 12516 15484
rect 11564 15262 11566 15314
rect 11618 15262 11620 15314
rect 9548 14140 9940 14196
rect 9548 12962 9604 14140
rect 9660 13972 9716 13982
rect 9660 13878 9716 13916
rect 9996 13860 10052 13870
rect 9996 13766 10052 13804
rect 11564 13858 11620 15262
rect 11900 15426 11956 15438
rect 11900 15374 11902 15426
rect 11954 15374 11956 15426
rect 11900 15204 11956 15374
rect 11900 15092 12292 15148
rect 12236 14530 12292 15092
rect 12460 15092 12516 15102
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 12236 14466 12292 14478
rect 12348 14532 12404 14542
rect 12348 14438 12404 14476
rect 12460 14530 12516 15036
rect 12460 14478 12462 14530
rect 12514 14478 12516 14530
rect 11564 13806 11566 13858
rect 11618 13806 11620 13858
rect 11564 13794 11620 13806
rect 12236 13858 12292 13870
rect 12236 13806 12238 13858
rect 12290 13806 12292 13858
rect 10332 13746 10388 13758
rect 10332 13694 10334 13746
rect 10386 13694 10388 13746
rect 10332 13636 10388 13694
rect 11452 13748 11508 13758
rect 11452 13654 11508 13692
rect 12012 13746 12068 13758
rect 12012 13694 12014 13746
rect 12066 13694 12068 13746
rect 10332 13570 10388 13580
rect 11004 13636 11060 13646
rect 9660 13188 9716 13198
rect 9660 13074 9716 13132
rect 9660 13022 9662 13074
rect 9714 13022 9716 13074
rect 9660 13010 9716 13022
rect 9548 12910 9550 12962
rect 9602 12910 9604 12962
rect 9548 12852 9604 12910
rect 9996 12962 10052 12974
rect 9996 12910 9998 12962
rect 10050 12910 10052 12962
rect 9548 12402 9604 12796
rect 9884 12850 9940 12862
rect 9884 12798 9886 12850
rect 9938 12798 9940 12850
rect 9884 12628 9940 12798
rect 9548 12350 9550 12402
rect 9602 12350 9604 12402
rect 9548 12338 9604 12350
rect 9772 12572 9884 12628
rect 9772 12402 9828 12572
rect 9884 12562 9940 12572
rect 9772 12350 9774 12402
rect 9826 12350 9828 12402
rect 9660 12068 9716 12078
rect 9660 11974 9716 12012
rect 9212 11396 9268 11452
rect 9212 11330 9268 11340
rect 9436 11394 9492 11452
rect 9436 11342 9438 11394
rect 9490 11342 9492 11394
rect 9436 11330 9492 11342
rect 9772 11394 9828 12350
rect 9996 12404 10052 12910
rect 10668 12962 10724 12974
rect 10668 12910 10670 12962
rect 10722 12910 10724 12962
rect 10444 12852 10500 12862
rect 10444 12758 10500 12796
rect 9996 12310 10052 12348
rect 10668 11956 10724 12910
rect 10668 11890 10724 11900
rect 10556 11508 10612 11518
rect 10556 11414 10612 11452
rect 9772 11342 9774 11394
rect 9826 11342 9828 11394
rect 9772 11330 9828 11342
rect 9100 11218 9156 11228
rect 10108 11284 10164 11294
rect 10164 11228 10276 11284
rect 10108 11190 10164 11228
rect 8764 10834 8932 10836
rect 8764 10782 8766 10834
rect 8818 10782 8932 10834
rect 8764 10780 8932 10782
rect 9660 11170 9716 11182
rect 9660 11118 9662 11170
rect 9714 11118 9716 11170
rect 8764 10770 8820 10780
rect 9660 10610 9716 11118
rect 9660 10558 9662 10610
rect 9714 10558 9716 10610
rect 9660 10546 9716 10558
rect 9772 11172 9828 11182
rect 9772 10610 9828 11116
rect 9772 10558 9774 10610
rect 9826 10558 9828 10610
rect 9772 10546 9828 10558
rect 9996 10724 10052 10734
rect 9996 10610 10052 10668
rect 9996 10558 9998 10610
rect 10050 10558 10052 10610
rect 9996 10546 10052 10558
rect 10108 10612 10164 10622
rect 10220 10612 10276 11228
rect 10556 10724 10612 10734
rect 10556 10630 10612 10668
rect 10332 10612 10388 10622
rect 10220 10556 10332 10612
rect 10108 10518 10164 10556
rect 10332 10546 10388 10556
rect 8876 10500 8932 10510
rect 8932 10444 9044 10500
rect 8876 10406 8932 10444
rect 8652 9998 8654 10050
rect 8706 9998 8708 10050
rect 8652 9986 8708 9998
rect 8988 9826 9044 10444
rect 8988 9774 8990 9826
rect 9042 9774 9044 9826
rect 8764 9602 8820 9614
rect 8764 9550 8766 9602
rect 8818 9550 8820 9602
rect 6300 8306 6356 8316
rect 8092 8372 8148 8382
rect 8764 8372 8820 9550
rect 8988 9604 9044 9774
rect 9436 9604 9492 9614
rect 8988 9602 9492 9604
rect 8988 9550 9438 9602
rect 9490 9550 9492 9602
rect 8988 9548 9492 9550
rect 9436 8708 9492 9548
rect 9436 8642 9492 8652
rect 10892 9042 10948 9054
rect 10892 8990 10894 9042
rect 10946 8990 10948 9042
rect 8876 8372 8932 8382
rect 8764 8370 8932 8372
rect 8764 8318 8878 8370
rect 8930 8318 8932 8370
rect 8764 8316 8932 8318
rect 8092 8258 8148 8316
rect 8876 8306 8932 8316
rect 10892 8372 10948 8990
rect 10892 8306 10948 8316
rect 11004 8370 11060 13580
rect 11340 13524 11396 13534
rect 11228 13468 11340 13524
rect 11228 12402 11284 13468
rect 11340 13458 11396 13468
rect 12012 13524 12068 13694
rect 12012 13458 12068 13468
rect 11788 12850 11844 12862
rect 11788 12798 11790 12850
rect 11842 12798 11844 12850
rect 11228 12350 11230 12402
rect 11282 12350 11284 12402
rect 11228 11732 11284 12350
rect 11564 12628 11620 12638
rect 11564 12402 11620 12572
rect 11564 12350 11566 12402
rect 11618 12350 11620 12402
rect 11564 12338 11620 12350
rect 11788 12404 11844 12798
rect 11900 12740 11956 12750
rect 11900 12646 11956 12684
rect 12236 12516 12292 13806
rect 12460 13748 12516 14478
rect 12460 13682 12516 13692
rect 12572 14530 12628 14542
rect 12572 14478 12574 14530
rect 12626 14478 12628 14530
rect 12572 12628 12628 14478
rect 12908 14530 12964 14542
rect 12908 14478 12910 14530
rect 12962 14478 12964 14530
rect 12908 14308 12964 14478
rect 12908 13746 12964 14252
rect 12908 13694 12910 13746
rect 12962 13694 12964 13746
rect 12908 13682 12964 13694
rect 12572 12562 12628 12572
rect 12236 12450 12292 12460
rect 11788 12338 11844 12348
rect 13132 12068 13188 19852
rect 13356 19842 13412 19852
rect 13468 20020 13524 20030
rect 13692 20020 13748 20030
rect 13468 20018 13748 20020
rect 13468 19966 13470 20018
rect 13522 19966 13694 20018
rect 13746 19966 13748 20018
rect 13468 19964 13748 19966
rect 13468 19460 13524 19964
rect 13692 19954 13748 19964
rect 13468 19394 13524 19404
rect 13580 19684 13636 19694
rect 13580 19346 13636 19628
rect 13580 19294 13582 19346
rect 13634 19294 13636 19346
rect 13580 19282 13636 19294
rect 13916 19460 13972 20078
rect 14476 20130 14532 20142
rect 14476 20078 14478 20130
rect 14530 20078 14532 20130
rect 14252 20020 14308 20030
rect 14252 19926 14308 19964
rect 14476 19908 14532 20078
rect 14588 20132 14644 20142
rect 14588 20038 14644 20076
rect 14476 19842 14532 19852
rect 14028 19796 14084 19806
rect 14028 19794 14420 19796
rect 14028 19742 14030 19794
rect 14082 19742 14420 19794
rect 14028 19740 14420 19742
rect 14028 19730 14084 19740
rect 14364 19572 14420 19740
rect 14364 19516 15092 19572
rect 13916 19404 14532 19460
rect 13916 18674 13972 19404
rect 14476 19346 14532 19404
rect 15036 19458 15092 19516
rect 15036 19406 15038 19458
rect 15090 19406 15092 19458
rect 15036 19394 15092 19406
rect 14476 19294 14478 19346
rect 14530 19294 14532 19346
rect 14476 19282 14532 19294
rect 14028 19236 14084 19246
rect 14028 19142 14084 19180
rect 14812 19234 14868 19246
rect 14812 19182 14814 19234
rect 14866 19182 14868 19234
rect 13916 18622 13918 18674
rect 13970 18622 13972 18674
rect 13916 18610 13972 18622
rect 13244 18562 13300 18574
rect 13244 18510 13246 18562
rect 13298 18510 13300 18562
rect 13244 18340 13300 18510
rect 14140 18562 14196 18574
rect 14140 18510 14142 18562
rect 14194 18510 14196 18562
rect 13692 18452 13748 18462
rect 13692 18358 13748 18396
rect 13244 18274 13300 18284
rect 14140 17892 14196 18510
rect 14252 18228 14308 18238
rect 14252 18134 14308 18172
rect 14812 17892 14868 19182
rect 15372 19236 15428 19246
rect 15372 19142 15428 19180
rect 14140 17836 14868 17892
rect 14476 17668 14532 17678
rect 13356 16770 13412 16782
rect 13356 16718 13358 16770
rect 13410 16718 13412 16770
rect 13356 13748 13412 16718
rect 13916 15540 13972 15550
rect 13692 15426 13748 15438
rect 13692 15374 13694 15426
rect 13746 15374 13748 15426
rect 13468 14420 13524 14430
rect 13468 14326 13524 14364
rect 13692 14308 13748 15374
rect 13916 15314 13972 15484
rect 14476 15426 14532 17612
rect 14476 15374 14478 15426
rect 14530 15374 14532 15426
rect 14476 15362 14532 15374
rect 13916 15262 13918 15314
rect 13970 15262 13972 15314
rect 13916 15250 13972 15262
rect 14364 15092 14420 15102
rect 14364 14998 14420 15036
rect 14588 14642 14644 17836
rect 16044 17668 16100 20638
rect 16380 20804 16436 20814
rect 16380 20690 16436 20748
rect 16380 20638 16382 20690
rect 16434 20638 16436 20690
rect 16380 20626 16436 20638
rect 16044 17602 16100 17612
rect 16828 18004 16884 18014
rect 16828 17666 16884 17948
rect 16828 17614 16830 17666
rect 16882 17614 16884 17666
rect 16828 17602 16884 17614
rect 16604 17554 16660 17566
rect 16604 17502 16606 17554
rect 16658 17502 16660 17554
rect 15484 17444 15540 17454
rect 15484 16994 15540 17388
rect 16492 17108 16548 17118
rect 16604 17108 16660 17502
rect 16716 17444 16772 17454
rect 16716 17350 16772 17388
rect 16492 17106 16660 17108
rect 16492 17054 16494 17106
rect 16546 17054 16660 17106
rect 16492 17052 16660 17054
rect 16492 17042 16548 17052
rect 15484 16942 15486 16994
rect 15538 16942 15540 16994
rect 15484 16930 15540 16942
rect 16716 16994 16772 17006
rect 16716 16942 16718 16994
rect 16770 16942 16772 16994
rect 16268 16884 16324 16894
rect 16268 16882 16548 16884
rect 16268 16830 16270 16882
rect 16322 16830 16548 16882
rect 16268 16828 16548 16830
rect 16268 16818 16324 16828
rect 16492 16210 16548 16828
rect 16716 16772 16772 16942
rect 16492 16158 16494 16210
rect 16546 16158 16548 16210
rect 16044 15540 16100 15550
rect 15372 15202 15428 15214
rect 15372 15150 15374 15202
rect 15426 15150 15428 15202
rect 14588 14590 14590 14642
rect 14642 14590 14644 14642
rect 14588 14578 14644 14590
rect 15036 14868 15092 14878
rect 14028 14532 14084 14542
rect 14476 14532 14532 14542
rect 14028 14438 14084 14476
rect 14140 14530 14532 14532
rect 14140 14478 14478 14530
rect 14530 14478 14532 14530
rect 14140 14476 14532 14478
rect 13692 14242 13748 14252
rect 13468 13972 13524 13982
rect 13468 13878 13524 13916
rect 13356 13682 13412 13692
rect 14028 13748 14084 13758
rect 14028 13654 14084 13692
rect 13804 13636 13860 13646
rect 13804 13542 13860 13580
rect 14140 13300 14196 14476
rect 14476 14466 14532 14476
rect 15036 14418 15092 14812
rect 15372 14868 15428 15150
rect 15372 14802 15428 14812
rect 16044 14754 16100 15484
rect 16380 15540 16436 15550
rect 16380 15446 16436 15484
rect 16492 15148 16548 16158
rect 16044 14702 16046 14754
rect 16098 14702 16100 14754
rect 16044 14690 16100 14702
rect 16268 15092 16548 15148
rect 16604 16716 16716 16772
rect 16604 15540 16660 16716
rect 16716 16706 16772 16716
rect 16828 16882 16884 16894
rect 16828 16830 16830 16882
rect 16882 16830 16884 16882
rect 16828 16324 16884 16830
rect 16828 16258 16884 16268
rect 16940 16322 16996 20860
rect 17276 20804 17332 20814
rect 17276 20710 17332 20748
rect 17164 20692 17220 20702
rect 17164 19124 17220 20636
rect 17388 20690 17444 21084
rect 17388 20638 17390 20690
rect 17442 20638 17444 20690
rect 17388 19348 17444 20638
rect 17388 19282 17444 19292
rect 17276 19124 17332 19134
rect 17612 19124 17668 22204
rect 18284 22194 18340 22206
rect 18508 22930 18564 22942
rect 18508 22878 18510 22930
rect 18562 22878 18564 22930
rect 17948 22148 18004 22158
rect 17836 22146 18004 22148
rect 17836 22094 17950 22146
rect 18002 22094 18004 22146
rect 17836 22092 18004 22094
rect 17164 19122 17444 19124
rect 17164 19070 17278 19122
rect 17330 19070 17444 19122
rect 17164 19068 17444 19070
rect 17276 19058 17332 19068
rect 17388 19012 17444 19068
rect 17388 18946 17444 18956
rect 17500 19122 17668 19124
rect 17500 19070 17614 19122
rect 17666 19070 17668 19122
rect 17500 19068 17668 19070
rect 17500 18788 17556 19068
rect 17612 19058 17668 19068
rect 17724 21028 17780 21038
rect 17164 18732 17556 18788
rect 17052 18452 17108 18462
rect 17052 17668 17108 18396
rect 17164 17890 17220 18732
rect 17164 17838 17166 17890
rect 17218 17838 17220 17890
rect 17164 17826 17220 17838
rect 17388 18340 17444 18350
rect 17164 17668 17220 17678
rect 17052 17666 17220 17668
rect 17052 17614 17166 17666
rect 17218 17614 17220 17666
rect 17052 17612 17220 17614
rect 16940 16270 16942 16322
rect 16994 16270 16996 16322
rect 15708 14532 15764 14542
rect 15484 14530 15764 14532
rect 15484 14478 15710 14530
rect 15762 14478 15764 14530
rect 15484 14476 15764 14478
rect 15036 14366 15038 14418
rect 15090 14366 15092 14418
rect 15036 14354 15092 14366
rect 15372 14420 15428 14430
rect 15372 14326 15428 14364
rect 15484 13970 15540 14476
rect 15708 14466 15764 14476
rect 16156 14420 16212 14430
rect 16156 14326 16212 14364
rect 15484 13918 15486 13970
rect 15538 13918 15540 13970
rect 15484 13906 15540 13918
rect 15596 14306 15652 14318
rect 15596 14254 15598 14306
rect 15650 14254 15652 14306
rect 15596 13972 15652 14254
rect 15596 13906 15652 13916
rect 14924 13748 14980 13758
rect 14700 13636 14756 13646
rect 14700 13542 14756 13580
rect 13692 13244 14196 13300
rect 14252 13524 14308 13534
rect 13580 12740 13636 12750
rect 13132 12002 13188 12012
rect 13468 12516 13524 12526
rect 11228 11666 11284 11676
rect 11900 11508 11956 11518
rect 11900 10836 11956 11452
rect 13468 11506 13524 12460
rect 13580 12404 13636 12684
rect 13580 12310 13636 12348
rect 13692 12402 13748 13244
rect 14252 13188 14308 13468
rect 13692 12350 13694 12402
rect 13746 12350 13748 12402
rect 13692 12338 13748 12350
rect 13804 13132 14308 13188
rect 13804 12402 13860 13132
rect 13804 12350 13806 12402
rect 13858 12350 13860 12402
rect 13804 12338 13860 12350
rect 13916 12850 13972 12862
rect 13916 12798 13918 12850
rect 13970 12798 13972 12850
rect 13916 11732 13972 12798
rect 14924 12404 14980 13692
rect 15036 13746 15092 13758
rect 15036 13694 15038 13746
rect 15090 13694 15092 13746
rect 15036 13524 15092 13694
rect 15596 13746 15652 13758
rect 15596 13694 15598 13746
rect 15650 13694 15652 13746
rect 15036 13458 15092 13468
rect 15260 13634 15316 13646
rect 15260 13582 15262 13634
rect 15314 13582 15316 13634
rect 14252 12402 14980 12404
rect 14252 12350 14926 12402
rect 14978 12350 14980 12402
rect 14252 12348 14980 12350
rect 14028 12292 14084 12302
rect 14028 12066 14084 12236
rect 14028 12014 14030 12066
rect 14082 12014 14084 12066
rect 14028 11956 14084 12014
rect 14028 11890 14084 11900
rect 14140 12180 14196 12190
rect 14028 11732 14084 11742
rect 13916 11676 14028 11732
rect 13468 11454 13470 11506
rect 13522 11454 13524 11506
rect 13468 11442 13524 11454
rect 12908 11396 12964 11406
rect 12348 10836 12404 10846
rect 11900 10834 12404 10836
rect 11900 10782 11902 10834
rect 11954 10782 12350 10834
rect 12402 10782 12404 10834
rect 11900 10780 12404 10782
rect 11900 10770 11956 10780
rect 12348 10770 12404 10780
rect 12124 10612 12180 10622
rect 12124 10518 12180 10556
rect 12572 10610 12628 10622
rect 12572 10558 12574 10610
rect 12626 10558 12628 10610
rect 12236 10498 12292 10510
rect 12236 10446 12238 10498
rect 12290 10446 12292 10498
rect 12124 9940 12180 9950
rect 12236 9940 12292 10446
rect 12572 10388 12628 10558
rect 12908 10610 12964 11340
rect 13580 11396 13636 11406
rect 13636 11340 13860 11396
rect 13580 11302 13636 11340
rect 12908 10558 12910 10610
rect 12962 10558 12964 10610
rect 12908 10546 12964 10558
rect 13356 10498 13412 10510
rect 13356 10446 13358 10498
rect 13410 10446 13412 10498
rect 13356 10388 13412 10446
rect 12572 10332 13412 10388
rect 12124 9938 12292 9940
rect 12124 9886 12126 9938
rect 12178 9886 12292 9938
rect 12124 9884 12292 9886
rect 12124 9874 12180 9884
rect 12012 9604 12068 9614
rect 11676 9602 12068 9604
rect 11676 9550 12014 9602
rect 12066 9550 12068 9602
rect 11676 9548 12068 9550
rect 11676 9154 11732 9548
rect 12012 9538 12068 9548
rect 11676 9102 11678 9154
rect 11730 9102 11732 9154
rect 11676 9090 11732 9102
rect 11004 8318 11006 8370
rect 11058 8318 11060 8370
rect 11004 8306 11060 8318
rect 11452 8372 11508 8382
rect 11452 8278 11508 8316
rect 13132 8372 13188 8382
rect 8092 8206 8094 8258
rect 8146 8206 8148 8258
rect 8092 8194 8148 8206
rect 13132 7476 13188 8316
rect 13132 7382 13188 7420
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 13356 6580 13412 10332
rect 13804 8930 13860 11340
rect 13804 8878 13806 8930
rect 13858 8878 13860 8930
rect 13804 8866 13860 8878
rect 14028 9938 14084 11676
rect 14140 11394 14196 12124
rect 14252 12178 14308 12348
rect 14924 12338 14980 12348
rect 15260 12404 15316 13582
rect 15484 13636 15540 13646
rect 15484 13542 15540 13580
rect 15596 12516 15652 13694
rect 15932 13748 15988 13758
rect 15932 13654 15988 13692
rect 15596 12450 15652 12460
rect 15260 12338 15316 12348
rect 15932 12290 15988 12302
rect 15932 12238 15934 12290
rect 15986 12238 15988 12290
rect 14252 12126 14254 12178
rect 14306 12126 14308 12178
rect 14252 12114 14308 12126
rect 14588 12178 14644 12190
rect 14588 12126 14590 12178
rect 14642 12126 14644 12178
rect 14588 12068 14644 12126
rect 15708 12180 15764 12190
rect 14588 12002 14644 12012
rect 15148 12068 15204 12078
rect 15148 11508 15204 12012
rect 15708 11844 15764 12124
rect 15708 11778 15764 11788
rect 15932 11508 15988 12238
rect 16268 12180 16324 15092
rect 16604 14084 16660 15484
rect 16828 15540 16884 15550
rect 16940 15540 16996 16270
rect 17052 16772 17108 16782
rect 17052 16210 17108 16716
rect 17052 16158 17054 16210
rect 17106 16158 17108 16210
rect 17052 16146 17108 16158
rect 16828 15538 16996 15540
rect 16828 15486 16830 15538
rect 16882 15486 16996 15538
rect 16828 15484 16996 15486
rect 16828 15474 16884 15484
rect 16716 15428 16772 15438
rect 16716 14754 16772 15372
rect 17164 15148 17220 17612
rect 17388 16996 17444 18284
rect 17612 18340 17668 18350
rect 17724 18340 17780 20972
rect 17836 20804 17892 22092
rect 17948 22082 18004 22092
rect 18396 21812 18452 21822
rect 17948 21700 18004 21710
rect 17948 21474 18004 21644
rect 18172 21588 18228 21598
rect 18172 21494 18228 21532
rect 17948 21422 17950 21474
rect 18002 21422 18004 21474
rect 17948 21028 18004 21422
rect 17948 20962 18004 20972
rect 18060 21364 18116 21374
rect 17836 20244 17892 20748
rect 18060 20802 18116 21308
rect 18060 20750 18062 20802
rect 18114 20750 18116 20802
rect 17948 20244 18004 20254
rect 17836 20242 18004 20244
rect 17836 20190 17950 20242
rect 18002 20190 18004 20242
rect 17836 20188 18004 20190
rect 17948 20178 18004 20188
rect 17836 20020 17892 20030
rect 18060 20020 18116 20750
rect 18396 21362 18452 21756
rect 18396 21310 18398 21362
rect 18450 21310 18452 21362
rect 18172 20692 18228 20702
rect 18172 20598 18228 20636
rect 18172 20244 18228 20254
rect 18172 20150 18228 20188
rect 18284 20020 18340 20030
rect 17836 20018 18116 20020
rect 17836 19966 17838 20018
rect 17890 19966 18116 20018
rect 17836 19964 18116 19966
rect 18172 19964 18284 20020
rect 17836 19954 17892 19964
rect 18060 19796 18116 19806
rect 17948 19740 18060 19796
rect 17836 18452 17892 18462
rect 17836 18358 17892 18396
rect 17668 18284 17780 18340
rect 17612 18274 17668 18284
rect 17836 17892 17892 17902
rect 17836 17798 17892 17836
rect 17724 16996 17780 17006
rect 17388 16994 17780 16996
rect 17388 16942 17726 16994
rect 17778 16942 17780 16994
rect 17388 16940 17780 16942
rect 17724 16930 17780 16940
rect 17948 16770 18004 19740
rect 18060 19730 18116 19740
rect 18060 19124 18116 19134
rect 18172 19124 18228 19964
rect 18284 19954 18340 19964
rect 18396 19236 18452 21310
rect 18508 19460 18564 22878
rect 18620 22484 18676 26236
rect 18620 22418 18676 22428
rect 18732 22260 18788 26348
rect 18732 21364 18788 22204
rect 18844 25506 18900 26460
rect 19180 26422 19236 26460
rect 18844 25454 18846 25506
rect 18898 25454 18900 25506
rect 18844 21588 18900 25454
rect 19068 26404 19124 26414
rect 18956 24052 19012 24062
rect 18956 23958 19012 23996
rect 19068 23268 19124 26348
rect 19292 26402 19348 27022
rect 19404 26740 19460 27692
rect 19404 26674 19460 26684
rect 19516 27074 19572 27086
rect 19516 27022 19518 27074
rect 19570 27022 19572 27074
rect 19516 26516 19572 27022
rect 19628 27076 19684 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19740 27076 19796 27086
rect 19628 27074 19796 27076
rect 19628 27022 19742 27074
rect 19794 27022 19796 27074
rect 19628 27020 19796 27022
rect 19740 27010 19796 27020
rect 20188 27074 20244 28364
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 20188 27010 20244 27022
rect 20412 27076 20468 27086
rect 20412 26982 20468 27020
rect 19628 26852 19684 26862
rect 19628 26758 19684 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19964 26516 20020 26526
rect 19292 26350 19294 26402
rect 19346 26350 19348 26402
rect 19292 26338 19348 26350
rect 19404 26514 20020 26516
rect 19404 26462 19966 26514
rect 20018 26462 20020 26514
rect 19404 26460 20020 26462
rect 19404 25508 19460 26460
rect 19964 26450 20020 26460
rect 19180 25452 19460 25508
rect 19180 25394 19236 25452
rect 19180 25342 19182 25394
rect 19234 25342 19236 25394
rect 19180 25330 19236 25342
rect 18956 23212 19124 23268
rect 18956 22930 19012 23212
rect 19068 23044 19124 23054
rect 19068 22950 19124 22988
rect 18956 22878 18958 22930
rect 19010 22878 19012 22930
rect 18956 22866 19012 22878
rect 19404 22708 19460 25452
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24164 20244 24174
rect 20188 24050 20244 24108
rect 20188 23998 20190 24050
rect 20242 23998 20244 24050
rect 20188 23986 20244 23998
rect 19852 23940 19908 23950
rect 19852 23846 19908 23884
rect 19628 23826 19684 23838
rect 19628 23774 19630 23826
rect 19682 23774 19684 23826
rect 19628 23604 19684 23774
rect 20188 23828 20244 23838
rect 20076 23716 20132 23754
rect 20188 23734 20244 23772
rect 20076 23650 20132 23660
rect 19628 23538 19684 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19516 23154 19572 23166
rect 19516 23102 19518 23154
rect 19570 23102 19572 23154
rect 19516 23044 19572 23102
rect 19516 22978 19572 22988
rect 19404 22652 19572 22708
rect 19404 22484 19460 22494
rect 19292 22148 19348 22158
rect 19180 22146 19348 22148
rect 19180 22094 19294 22146
rect 19346 22094 19348 22146
rect 19180 22092 19348 22094
rect 19180 21588 19236 22092
rect 19292 22082 19348 22092
rect 19292 21700 19348 21710
rect 19292 21606 19348 21644
rect 18844 21532 19012 21588
rect 18844 21364 18900 21374
rect 18732 21362 18900 21364
rect 18732 21310 18846 21362
rect 18898 21310 18900 21362
rect 18732 21308 18900 21310
rect 18844 21298 18900 21308
rect 18844 20916 18900 20926
rect 18844 20822 18900 20860
rect 18620 20580 18676 20590
rect 18620 20486 18676 20524
rect 18956 20132 19012 21532
rect 19180 21522 19236 21532
rect 19404 21474 19460 22428
rect 19404 21422 19406 21474
rect 19458 21422 19460 21474
rect 19404 21410 19460 21422
rect 19068 21364 19124 21374
rect 19068 21270 19124 21308
rect 19516 21028 19572 22652
rect 19628 22372 19684 22382
rect 19628 22278 19684 22316
rect 20524 22372 20580 32060
rect 20748 31892 20804 31902
rect 20748 29538 20804 31836
rect 21420 31780 21476 31790
rect 21420 31666 21476 31724
rect 22428 31780 22484 33070
rect 22428 31714 22484 31724
rect 21420 31614 21422 31666
rect 21474 31614 21476 31666
rect 21420 31602 21476 31614
rect 21532 31666 21588 31678
rect 21532 31614 21534 31666
rect 21586 31614 21588 31666
rect 20860 31554 20916 31566
rect 20860 31502 20862 31554
rect 20914 31502 20916 31554
rect 20860 30100 20916 31502
rect 21196 31556 21252 31566
rect 21532 31556 21588 31614
rect 21196 31554 21364 31556
rect 21196 31502 21198 31554
rect 21250 31502 21364 31554
rect 21196 31500 21364 31502
rect 21196 31490 21252 31500
rect 20860 30006 20916 30044
rect 21196 29540 21252 29550
rect 20748 29486 20750 29538
rect 20802 29486 20804 29538
rect 20748 29474 20804 29486
rect 20860 29538 21252 29540
rect 20860 29486 21198 29538
rect 21250 29486 21252 29538
rect 20860 29484 21252 29486
rect 20860 29426 20916 29484
rect 21196 29474 21252 29484
rect 20860 29374 20862 29426
rect 20914 29374 20916 29426
rect 20860 29362 20916 29374
rect 21084 29316 21140 29326
rect 20636 27074 20692 27086
rect 20636 27022 20638 27074
rect 20690 27022 20692 27074
rect 20636 26180 20692 27022
rect 20748 26964 20804 27002
rect 20748 26898 20804 26908
rect 20972 26180 21028 26190
rect 20636 26178 21028 26180
rect 20636 26126 20974 26178
rect 21026 26126 21028 26178
rect 20636 26124 21028 26126
rect 20860 24610 20916 26124
rect 20972 26114 21028 26124
rect 20860 24558 20862 24610
rect 20914 24558 20916 24610
rect 20636 24388 20692 24398
rect 20636 23826 20692 24332
rect 20748 24164 20804 24174
rect 20748 24050 20804 24108
rect 20748 23998 20750 24050
rect 20802 23998 20804 24050
rect 20748 23986 20804 23998
rect 20636 23774 20638 23826
rect 20690 23774 20692 23826
rect 20636 23762 20692 23774
rect 20524 22306 20580 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20860 21700 20916 24558
rect 20748 21644 20916 21700
rect 20972 22372 21028 22382
rect 20748 21476 20804 21644
rect 18956 20066 19012 20076
rect 19180 20972 19572 21028
rect 20524 21420 20804 21476
rect 20860 21476 20916 21486
rect 20972 21476 21028 22316
rect 20860 21474 21028 21476
rect 20860 21422 20862 21474
rect 20914 21422 21028 21474
rect 20860 21420 21028 21422
rect 18956 19908 19012 19918
rect 19068 19908 19124 19918
rect 18956 19906 19068 19908
rect 18956 19854 18958 19906
rect 19010 19854 19068 19906
rect 18956 19852 19068 19854
rect 18956 19842 19012 19852
rect 18508 19404 18676 19460
rect 18508 19236 18564 19246
rect 18396 19234 18564 19236
rect 18396 19182 18510 19234
rect 18562 19182 18564 19234
rect 18396 19180 18564 19182
rect 18508 19170 18564 19180
rect 18060 19122 18228 19124
rect 18060 19070 18062 19122
rect 18114 19070 18228 19122
rect 18060 19068 18228 19070
rect 18060 19058 18116 19068
rect 18620 18788 18676 19404
rect 18956 19234 19012 19246
rect 18956 19182 18958 19234
rect 19010 19182 19012 19234
rect 18956 19012 19012 19182
rect 18956 18946 19012 18956
rect 18396 18732 18676 18788
rect 18284 18452 18340 18462
rect 18396 18452 18452 18732
rect 18284 18450 18452 18452
rect 18284 18398 18286 18450
rect 18338 18398 18452 18450
rect 18284 18396 18452 18398
rect 18508 18564 18564 18574
rect 18284 18386 18340 18396
rect 18396 18226 18452 18238
rect 18396 18174 18398 18226
rect 18450 18174 18452 18226
rect 18396 17666 18452 18174
rect 18396 17614 18398 17666
rect 18450 17614 18452 17666
rect 18396 17602 18452 17614
rect 18284 17556 18340 17566
rect 17948 16718 17950 16770
rect 18002 16718 18004 16770
rect 17948 16706 18004 16718
rect 18060 17554 18340 17556
rect 18060 17502 18286 17554
rect 18338 17502 18340 17554
rect 18060 17500 18340 17502
rect 17612 16322 17668 16334
rect 17612 16270 17614 16322
rect 17666 16270 17668 16322
rect 17612 16210 17668 16270
rect 17948 16324 18004 16334
rect 18060 16324 18116 17500
rect 18284 17490 18340 17500
rect 18004 16268 18116 16324
rect 18172 16658 18228 16670
rect 18172 16606 18174 16658
rect 18226 16606 18228 16658
rect 17948 16230 18004 16268
rect 17612 16158 17614 16210
rect 17666 16158 17668 16210
rect 17612 15876 17668 16158
rect 18172 16100 18228 16606
rect 17164 15092 17332 15148
rect 16716 14702 16718 14754
rect 16770 14702 16772 14754
rect 16716 14690 16772 14702
rect 16828 14420 16884 14430
rect 16828 14418 17108 14420
rect 16828 14366 16830 14418
rect 16882 14366 17108 14418
rect 16828 14364 17108 14366
rect 16828 14354 16884 14364
rect 16716 14308 16772 14318
rect 16716 14214 16772 14252
rect 16604 14028 16996 14084
rect 16604 13972 16660 14028
rect 16380 13916 16660 13972
rect 16380 13858 16436 13916
rect 16380 13806 16382 13858
rect 16434 13806 16436 13858
rect 16380 13794 16436 13806
rect 16828 13858 16884 13870
rect 16828 13806 16830 13858
rect 16882 13806 16884 13858
rect 16604 13746 16660 13758
rect 16604 13694 16606 13746
rect 16658 13694 16660 13746
rect 16156 12124 16324 12180
rect 16380 12292 16436 12302
rect 16604 12292 16660 13694
rect 16828 13748 16884 13806
rect 16828 13682 16884 13692
rect 16716 13634 16772 13646
rect 16716 13582 16718 13634
rect 16770 13582 16772 13634
rect 16716 12964 16772 13582
rect 16716 12898 16772 12908
rect 16380 12290 16660 12292
rect 16380 12238 16382 12290
rect 16434 12238 16660 12290
rect 16380 12236 16660 12238
rect 16156 11732 16212 12124
rect 16156 11666 16212 11676
rect 16380 11508 16436 12236
rect 16492 12066 16548 12078
rect 16492 12014 16494 12066
rect 16546 12014 16548 12066
rect 16492 11620 16548 12014
rect 16604 12068 16660 12078
rect 16604 11974 16660 12012
rect 16940 11732 16996 14028
rect 17052 13412 17108 14364
rect 17164 13412 17220 13422
rect 17052 13356 17164 13412
rect 17164 13346 17220 13356
rect 17276 12292 17332 15092
rect 17388 14980 17444 14990
rect 17388 14418 17444 14924
rect 17612 14532 17668 15820
rect 17948 16044 18228 16100
rect 18396 16658 18452 16670
rect 18396 16606 18398 16658
rect 18450 16606 18452 16658
rect 17948 15538 18004 16044
rect 18284 15986 18340 15998
rect 18284 15934 18286 15986
rect 18338 15934 18340 15986
rect 18060 15876 18116 15886
rect 18060 15782 18116 15820
rect 17948 15486 17950 15538
rect 18002 15486 18004 15538
rect 17724 15426 17780 15438
rect 17724 15374 17726 15426
rect 17778 15374 17780 15426
rect 17724 14644 17780 15374
rect 17948 14756 18004 15486
rect 18172 15428 18228 15438
rect 18172 15334 18228 15372
rect 18060 15092 18116 15102
rect 18060 14998 18116 15036
rect 17948 14690 18004 14700
rect 17836 14644 17892 14654
rect 17724 14642 17892 14644
rect 17724 14590 17838 14642
rect 17890 14590 17892 14642
rect 17724 14588 17892 14590
rect 17836 14578 17892 14588
rect 17612 14476 17780 14532
rect 17388 14366 17390 14418
rect 17442 14366 17444 14418
rect 17388 13860 17444 14366
rect 17388 13794 17444 13804
rect 17500 14308 17556 14318
rect 16940 11666 16996 11676
rect 17052 12236 17332 12292
rect 17500 12292 17556 14252
rect 17612 14306 17668 14318
rect 17612 14254 17614 14306
rect 17666 14254 17668 14306
rect 17612 13748 17668 14254
rect 17724 14308 17780 14476
rect 17948 14420 18004 14430
rect 18004 14364 18228 14420
rect 17948 14326 18004 14364
rect 17836 14308 17892 14318
rect 17724 14306 17892 14308
rect 17724 14254 17838 14306
rect 17890 14254 17892 14306
rect 17724 14252 17892 14254
rect 17836 13860 17892 14252
rect 17836 13794 17892 13804
rect 17948 13860 18004 13870
rect 17948 13858 18116 13860
rect 17948 13806 17950 13858
rect 18002 13806 18116 13858
rect 17948 13804 18116 13806
rect 17948 13794 18004 13804
rect 17612 13682 17668 13692
rect 17724 13746 17780 13758
rect 17724 13694 17726 13746
rect 17778 13694 17780 13746
rect 17612 12292 17668 12302
rect 17500 12290 17668 12292
rect 17500 12238 17614 12290
rect 17666 12238 17668 12290
rect 17500 12236 17668 12238
rect 16492 11554 16548 11564
rect 15932 11452 16436 11508
rect 15148 11414 15204 11452
rect 14140 11342 14142 11394
rect 14194 11342 14196 11394
rect 14140 11330 14196 11342
rect 16380 11396 16436 11452
rect 16828 11396 16884 11406
rect 16380 11340 16828 11396
rect 16828 11302 16884 11340
rect 14588 11284 14644 11294
rect 16940 11284 16996 11294
rect 14644 11228 14756 11284
rect 14588 11218 14644 11228
rect 14028 9886 14030 9938
rect 14082 9886 14084 9938
rect 13916 8372 13972 8382
rect 14028 8372 14084 9886
rect 14252 8932 14308 8942
rect 14252 8930 14644 8932
rect 14252 8878 14254 8930
rect 14306 8878 14644 8930
rect 14252 8876 14644 8878
rect 14252 8866 14308 8876
rect 14364 8708 14420 8718
rect 14252 8372 14308 8382
rect 13972 8316 14084 8372
rect 14140 8370 14308 8372
rect 14140 8318 14254 8370
rect 14306 8318 14308 8370
rect 14140 8316 14308 8318
rect 13916 8306 13972 8316
rect 14028 8148 14084 8158
rect 14028 8054 14084 8092
rect 13916 7588 13972 7598
rect 14140 7588 14196 8316
rect 14252 8306 14308 8316
rect 14364 8034 14420 8652
rect 14588 8482 14644 8876
rect 14588 8430 14590 8482
rect 14642 8430 14644 8482
rect 14588 8418 14644 8430
rect 14700 8930 14756 11228
rect 16940 11190 16996 11228
rect 16044 11172 16100 11182
rect 16044 9938 16100 11116
rect 17052 10724 17108 12236
rect 17612 12226 17668 12236
rect 17388 12180 17444 12190
rect 17164 12178 17444 12180
rect 17164 12126 17390 12178
rect 17442 12126 17444 12178
rect 17164 12124 17444 12126
rect 17164 11394 17220 12124
rect 17388 12114 17444 12124
rect 17164 11342 17166 11394
rect 17218 11342 17220 11394
rect 17164 11330 17220 11342
rect 17500 12066 17556 12078
rect 17500 12014 17502 12066
rect 17554 12014 17556 12066
rect 17388 11172 17444 11182
rect 17388 11078 17444 11116
rect 17052 10658 17108 10668
rect 17500 10276 17556 12014
rect 17724 11844 17780 13694
rect 18060 13412 18116 13804
rect 18172 13858 18228 14364
rect 18284 13972 18340 15934
rect 18396 15428 18452 16606
rect 18508 16548 18564 18508
rect 18620 18004 18676 18732
rect 18844 18676 18900 18686
rect 19068 18676 19124 19852
rect 18900 18620 19124 18676
rect 18844 18226 18900 18620
rect 18844 18174 18846 18226
rect 18898 18174 18900 18226
rect 18844 18162 18900 18174
rect 18620 17938 18676 17948
rect 19068 17892 19124 17902
rect 19068 17798 19124 17836
rect 18508 16482 18564 16492
rect 18620 17666 18676 17678
rect 18620 17614 18622 17666
rect 18674 17614 18676 17666
rect 18620 17556 18676 17614
rect 18956 17556 19012 17566
rect 18620 17554 19012 17556
rect 18620 17502 18958 17554
rect 19010 17502 19012 17554
rect 18620 17500 19012 17502
rect 18396 15362 18452 15372
rect 18508 16324 18564 16334
rect 18508 15314 18564 16268
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 15250 18564 15262
rect 18508 14980 18564 14990
rect 18620 14980 18676 17500
rect 18956 17490 19012 17500
rect 19180 16996 19236 20972
rect 20076 20802 20132 20814
rect 20076 20750 20078 20802
rect 20130 20750 20132 20802
rect 19516 20690 19572 20702
rect 19740 20692 19796 20702
rect 19516 20638 19518 20690
rect 19570 20638 19572 20690
rect 19292 20132 19348 20142
rect 19292 20038 19348 20076
rect 19516 19348 19572 20638
rect 19628 20690 19796 20692
rect 19628 20638 19742 20690
rect 19794 20638 19796 20690
rect 19628 20636 19796 20638
rect 19628 20244 19684 20636
rect 19740 20626 19796 20636
rect 20076 20580 20132 20750
rect 20076 20524 20244 20580
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19628 20188 19796 20244
rect 19740 20132 19796 20188
rect 19740 20066 19796 20076
rect 19628 20018 19684 20030
rect 19628 19966 19630 20018
rect 19682 19966 19684 20018
rect 19628 19908 19684 19966
rect 19628 19842 19684 19852
rect 20188 20018 20244 20524
rect 20412 20132 20468 20142
rect 20412 20038 20468 20076
rect 20188 19966 20190 20018
rect 20242 19966 20244 20018
rect 20188 19348 20244 19966
rect 19516 19292 19684 19348
rect 20188 19292 20468 19348
rect 19516 19122 19572 19134
rect 19516 19070 19518 19122
rect 19570 19070 19572 19122
rect 19404 19012 19460 19022
rect 19404 18918 19460 18956
rect 19404 18116 19460 18126
rect 19068 16940 19236 16996
rect 19292 18004 19348 18014
rect 19068 16772 19124 16940
rect 19068 16706 19124 16716
rect 19292 16772 19348 17948
rect 19404 17556 19460 18060
rect 19516 17778 19572 19070
rect 19628 19124 19684 19292
rect 19628 19058 19684 19068
rect 19964 19234 20020 19246
rect 19964 19182 19966 19234
rect 20018 19182 20020 19234
rect 19964 19124 20020 19182
rect 19964 19058 20020 19068
rect 20188 19122 20244 19134
rect 20188 19070 20190 19122
rect 20242 19070 20244 19122
rect 20188 18900 20244 19070
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20188 18834 20244 18844
rect 20300 19122 20356 19134
rect 20300 19070 20302 19122
rect 20354 19070 20356 19122
rect 20300 19012 20356 19070
rect 19836 18778 20100 18788
rect 20076 18676 20132 18686
rect 20300 18676 20356 18956
rect 20076 18674 20356 18676
rect 20076 18622 20078 18674
rect 20130 18622 20356 18674
rect 20076 18620 20356 18622
rect 20076 18610 20132 18620
rect 19740 18564 19796 18574
rect 19740 18470 19796 18508
rect 20412 18564 20468 19292
rect 20412 18498 20468 18508
rect 20524 18452 20580 21420
rect 20636 20580 20692 20590
rect 20636 20018 20692 20524
rect 20636 19966 20638 20018
rect 20690 19966 20692 20018
rect 20636 19954 20692 19966
rect 20748 20244 20804 20254
rect 20748 20018 20804 20188
rect 20748 19966 20750 20018
rect 20802 19966 20804 20018
rect 20748 19954 20804 19966
rect 20860 20020 20916 21420
rect 20972 20242 21028 20254
rect 20972 20190 20974 20242
rect 21026 20190 21028 20242
rect 20972 20132 21028 20190
rect 20972 20066 21028 20076
rect 20860 19954 20916 19964
rect 21084 19796 21140 29260
rect 21308 29204 21364 31500
rect 21532 31490 21588 31500
rect 21868 31554 21924 31566
rect 21868 31502 21870 31554
rect 21922 31502 21924 31554
rect 21868 30100 21924 31502
rect 22204 31554 22260 31566
rect 22204 31502 22206 31554
rect 22258 31502 22260 31554
rect 22204 31220 22260 31502
rect 22204 31154 22260 31164
rect 21532 29988 21588 29998
rect 21420 29428 21476 29438
rect 21420 29334 21476 29372
rect 21308 29148 21476 29204
rect 21308 27188 21364 27198
rect 21196 24724 21252 24734
rect 21196 24630 21252 24668
rect 21308 23492 21364 27132
rect 21420 23940 21476 29148
rect 21532 25284 21588 29932
rect 21868 29986 21924 30044
rect 22204 30324 22260 30334
rect 22204 30098 22260 30268
rect 22204 30046 22206 30098
rect 22258 30046 22260 30098
rect 22204 30034 22260 30046
rect 21868 29934 21870 29986
rect 21922 29934 21924 29986
rect 21532 25218 21588 25228
rect 21756 29426 21812 29438
rect 21756 29374 21758 29426
rect 21810 29374 21812 29426
rect 21420 23874 21476 23884
rect 21308 23426 21364 23436
rect 21644 23716 21700 23726
rect 21308 23268 21364 23278
rect 21308 22260 21364 23212
rect 21644 22370 21700 23660
rect 21644 22318 21646 22370
rect 21698 22318 21700 22370
rect 21644 22306 21700 22318
rect 21308 22258 21476 22260
rect 21308 22206 21310 22258
rect 21362 22206 21476 22258
rect 21308 22204 21476 22206
rect 21308 22194 21364 22204
rect 21308 20804 21364 20814
rect 21196 20802 21364 20804
rect 21196 20750 21310 20802
rect 21362 20750 21364 20802
rect 21196 20748 21364 20750
rect 21196 20580 21252 20748
rect 21308 20738 21364 20748
rect 21196 20018 21252 20524
rect 21420 20132 21476 22204
rect 21532 21476 21588 21486
rect 21532 21026 21588 21420
rect 21756 21252 21812 29374
rect 21868 29316 21924 29934
rect 22540 29428 22596 36204
rect 23324 35922 23380 36316
rect 23324 35870 23326 35922
rect 23378 35870 23380 35922
rect 23324 35858 23380 35870
rect 22988 35588 23044 35598
rect 22988 32676 23044 35532
rect 23100 34916 23156 34926
rect 23436 34916 23492 36988
rect 24668 36372 24724 37886
rect 25116 37940 25172 37950
rect 25116 37846 25172 37884
rect 24892 37826 24948 37838
rect 24892 37774 24894 37826
rect 24946 37774 24948 37826
rect 24892 36594 24948 37774
rect 25340 37156 25396 37998
rect 26124 38050 26180 38062
rect 26124 37998 26126 38050
rect 26178 37998 26180 38050
rect 25564 37156 25620 37166
rect 25676 37156 25732 37166
rect 25340 37154 25676 37156
rect 25340 37102 25566 37154
rect 25618 37102 25676 37154
rect 25340 37100 25676 37102
rect 25564 37090 25620 37100
rect 24892 36542 24894 36594
rect 24946 36542 24948 36594
rect 24892 36530 24948 36542
rect 24668 36306 24724 36316
rect 25452 36482 25508 36494
rect 25452 36430 25454 36482
rect 25506 36430 25508 36482
rect 23548 35698 23604 35710
rect 23548 35646 23550 35698
rect 23602 35646 23604 35698
rect 23548 35588 23604 35646
rect 23548 35522 23604 35532
rect 24780 35588 24836 35598
rect 24780 35494 24836 35532
rect 23100 34914 23492 34916
rect 23100 34862 23102 34914
rect 23154 34862 23492 34914
rect 23100 34860 23492 34862
rect 23100 33460 23156 34860
rect 23772 34804 23828 34814
rect 23772 34802 23940 34804
rect 23772 34750 23774 34802
rect 23826 34750 23940 34802
rect 23772 34748 23940 34750
rect 23772 34738 23828 34748
rect 23436 34692 23492 34702
rect 23436 34354 23492 34636
rect 23436 34302 23438 34354
rect 23490 34302 23492 34354
rect 23436 34132 23492 34302
rect 23884 34354 23940 34748
rect 23884 34302 23886 34354
rect 23938 34302 23940 34354
rect 23884 34290 23940 34302
rect 23660 34132 23716 34142
rect 24108 34132 24164 34142
rect 23436 34130 24052 34132
rect 23436 34078 23662 34130
rect 23714 34078 24052 34130
rect 23436 34076 24052 34078
rect 23660 34066 23716 34076
rect 23100 33394 23156 33404
rect 22988 31220 23044 32620
rect 23212 32788 23268 32798
rect 23212 31778 23268 32732
rect 23996 32788 24052 34076
rect 24108 34038 24164 34076
rect 24332 34132 24388 34142
rect 25452 34132 25508 36430
rect 25676 34244 25732 37100
rect 26124 36932 26180 37998
rect 26572 38050 26628 38108
rect 26572 37998 26574 38050
rect 26626 37998 26628 38050
rect 26572 37940 26628 37998
rect 26572 37874 26628 37884
rect 26684 37938 26740 37950
rect 26684 37886 26686 37938
rect 26738 37886 26740 37938
rect 26684 37604 26740 37886
rect 26460 37548 26740 37604
rect 26460 37268 26516 37548
rect 26124 36866 26180 36876
rect 26236 37266 26516 37268
rect 26236 37214 26462 37266
rect 26514 37214 26516 37266
rect 26236 37212 26516 37214
rect 25788 36596 25844 36606
rect 26236 36596 26292 37212
rect 26460 37202 26516 37212
rect 26572 37378 26628 37390
rect 26572 37326 26574 37378
rect 26626 37326 26628 37378
rect 25788 36594 26292 36596
rect 25788 36542 25790 36594
rect 25842 36542 26292 36594
rect 25788 36540 26292 36542
rect 26460 36932 26516 36942
rect 26460 36596 26516 36876
rect 25788 36530 25844 36540
rect 26460 36502 26516 36540
rect 25788 35364 25844 35374
rect 25788 34468 25844 35308
rect 26572 35140 26628 37326
rect 26684 36484 26740 36494
rect 26796 36484 26852 38108
rect 27356 37940 27412 37950
rect 27356 37846 27412 37884
rect 27468 37490 27524 38612
rect 28028 38162 28084 39452
rect 29148 39394 29204 39406
rect 29148 39342 29150 39394
rect 29202 39342 29204 39394
rect 28252 38836 28308 38846
rect 28252 38742 28308 38780
rect 28812 38724 28868 38734
rect 28028 38110 28030 38162
rect 28082 38110 28084 38162
rect 28028 38098 28084 38110
rect 28364 38722 28868 38724
rect 28364 38670 28814 38722
rect 28866 38670 28868 38722
rect 28364 38668 28868 38670
rect 27468 37438 27470 37490
rect 27522 37438 27524 37490
rect 27468 37426 27524 37438
rect 27916 38052 27972 38062
rect 27916 37492 27972 37996
rect 28364 38050 28420 38668
rect 28812 38658 28868 38668
rect 28364 37998 28366 38050
rect 28418 37998 28420 38050
rect 28364 37986 28420 37998
rect 28588 37940 28644 37950
rect 28140 37828 28196 37838
rect 28140 37734 28196 37772
rect 28028 37492 28084 37502
rect 27916 37490 28084 37492
rect 27916 37438 28030 37490
rect 28082 37438 28084 37490
rect 27916 37436 28084 37438
rect 27356 37268 27412 37278
rect 27020 37266 27412 37268
rect 27020 37214 27358 37266
rect 27410 37214 27412 37266
rect 27020 37212 27412 37214
rect 27020 36706 27076 37212
rect 27356 37202 27412 37212
rect 27916 37156 27972 37436
rect 28028 37426 28084 37436
rect 27916 37090 27972 37100
rect 27020 36654 27022 36706
rect 27074 36654 27076 36706
rect 27020 36642 27076 36654
rect 26684 36482 26852 36484
rect 26684 36430 26686 36482
rect 26738 36430 26852 36482
rect 26684 36428 26852 36430
rect 26684 35252 26740 36428
rect 27244 36260 27300 36270
rect 26796 35698 26852 35710
rect 26796 35646 26798 35698
rect 26850 35646 26852 35698
rect 26796 35588 26852 35646
rect 26796 35522 26852 35532
rect 26908 35588 26964 35598
rect 26684 35186 26740 35196
rect 25900 35084 26628 35140
rect 25900 35026 25956 35084
rect 25900 34974 25902 35026
rect 25954 34974 25956 35026
rect 25900 34962 25956 34974
rect 26236 34914 26292 34926
rect 26236 34862 26238 34914
rect 26290 34862 26292 34914
rect 25788 34412 26068 34468
rect 25788 34244 25844 34254
rect 25676 34242 25956 34244
rect 25676 34190 25790 34242
rect 25842 34190 25956 34242
rect 25676 34188 25956 34190
rect 25788 34178 25844 34188
rect 24332 34130 24500 34132
rect 24332 34078 24334 34130
rect 24386 34078 24500 34130
rect 24332 34076 24500 34078
rect 24332 34066 24388 34076
rect 23996 32786 24388 32788
rect 23996 32734 23998 32786
rect 24050 32734 24388 32786
rect 23996 32732 24388 32734
rect 23996 32722 24052 32732
rect 24332 32674 24388 32732
rect 24332 32622 24334 32674
rect 24386 32622 24388 32674
rect 24332 32610 24388 32622
rect 23548 31892 23604 31902
rect 23212 31726 23214 31778
rect 23266 31726 23268 31778
rect 23212 31714 23268 31726
rect 23324 31780 23380 31790
rect 22988 31154 23044 31164
rect 22988 30324 23044 30334
rect 22988 30230 23044 30268
rect 22764 30210 22820 30222
rect 22764 30158 22766 30210
rect 22818 30158 22820 30210
rect 22764 29988 22820 30158
rect 23324 30210 23380 31724
rect 23548 31778 23604 31836
rect 23548 31726 23550 31778
rect 23602 31726 23604 31778
rect 23548 31714 23604 31726
rect 24108 31780 24164 31790
rect 24108 31686 24164 31724
rect 23772 31666 23828 31678
rect 23772 31614 23774 31666
rect 23826 31614 23828 31666
rect 23548 31556 23604 31566
rect 23548 31462 23604 31500
rect 23772 30884 23828 31614
rect 23884 31556 23940 31566
rect 23884 30996 23940 31500
rect 24332 30996 24388 31006
rect 23884 30994 24164 30996
rect 23884 30942 23886 30994
rect 23938 30942 24164 30994
rect 23884 30940 24164 30942
rect 23884 30930 23940 30940
rect 23772 30818 23828 30828
rect 23324 30158 23326 30210
rect 23378 30158 23380 30210
rect 23324 30146 23380 30158
rect 24108 30324 24164 30940
rect 24332 30902 24388 30940
rect 22764 29922 22820 29932
rect 23324 29540 23380 29550
rect 22764 29428 22820 29438
rect 22540 29426 22820 29428
rect 22540 29374 22766 29426
rect 22818 29374 22820 29426
rect 22540 29372 22820 29374
rect 21868 29250 21924 29260
rect 22428 28420 22484 28430
rect 22764 28420 22820 29372
rect 23324 29426 23380 29484
rect 23324 29374 23326 29426
rect 23378 29374 23380 29426
rect 23324 29362 23380 29374
rect 24108 29426 24164 30268
rect 24108 29374 24110 29426
rect 24162 29374 24164 29426
rect 24108 29362 24164 29374
rect 23772 29314 23828 29326
rect 23772 29262 23774 29314
rect 23826 29262 23828 29314
rect 22428 28418 22820 28420
rect 22428 28366 22430 28418
rect 22482 28366 22820 28418
rect 22428 28364 22820 28366
rect 23660 28642 23716 28654
rect 23660 28590 23662 28642
rect 23714 28590 23716 28642
rect 23660 28420 23716 28590
rect 22428 28354 22484 28364
rect 22540 27970 22596 28364
rect 22540 27918 22542 27970
rect 22594 27918 22596 27970
rect 22540 27300 22596 27918
rect 22540 27234 22596 27244
rect 22876 27858 22932 27870
rect 22876 27806 22878 27858
rect 22930 27806 22932 27858
rect 22876 26908 22932 27806
rect 23324 27860 23380 27870
rect 22876 26852 23268 26908
rect 23212 26290 23268 26852
rect 23212 26238 23214 26290
rect 23266 26238 23268 26290
rect 22764 25396 22820 25406
rect 22764 25302 22820 25340
rect 23212 25396 23268 26238
rect 23212 25330 23268 25340
rect 22428 25282 22484 25294
rect 22428 25230 22430 25282
rect 22482 25230 22484 25282
rect 22428 25060 22484 25230
rect 22204 25004 22484 25060
rect 22092 24724 22148 24734
rect 22204 24724 22260 25004
rect 22316 24836 22372 24846
rect 22316 24742 22372 24780
rect 22148 24668 22260 24724
rect 22092 23940 22148 24668
rect 22316 23940 22372 23950
rect 22092 23938 22372 23940
rect 22092 23886 22318 23938
rect 22370 23886 22372 23938
rect 22092 23884 22372 23886
rect 21868 23714 21924 23726
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21868 23380 21924 23662
rect 21868 23314 21924 23324
rect 22092 23714 22148 23726
rect 22092 23662 22094 23714
rect 22146 23662 22148 23714
rect 22092 23156 22148 23662
rect 22316 23716 22372 23884
rect 23100 23940 23156 23950
rect 23100 23846 23156 23884
rect 22316 23650 22372 23660
rect 22764 23828 22820 23838
rect 22764 23380 22820 23772
rect 22876 23716 22932 23726
rect 22876 23714 23156 23716
rect 22876 23662 22878 23714
rect 22930 23662 23156 23714
rect 22876 23660 23156 23662
rect 22876 23650 22932 23660
rect 23100 23380 23156 23660
rect 22764 23324 23044 23380
rect 22092 21924 22148 23100
rect 22988 22482 23044 23324
rect 23100 23314 23156 23324
rect 23324 23268 23380 27804
rect 23548 27076 23604 27086
rect 23436 26964 23492 27002
rect 23436 26898 23492 26908
rect 23548 26514 23604 27020
rect 23548 26462 23550 26514
rect 23602 26462 23604 26514
rect 23548 26450 23604 26462
rect 23660 24948 23716 28364
rect 23772 27412 23828 29262
rect 24220 28756 24276 28766
rect 24444 28756 24500 34076
rect 25116 33460 25172 33470
rect 25116 33346 25172 33404
rect 25116 33294 25118 33346
rect 25170 33294 25172 33346
rect 25116 33282 25172 33294
rect 24556 32674 24612 32686
rect 24556 32622 24558 32674
rect 24610 32622 24612 32674
rect 24556 30324 24612 32622
rect 24668 32452 24724 32462
rect 24668 32358 24724 32396
rect 24668 31778 24724 31790
rect 24668 31726 24670 31778
rect 24722 31726 24724 31778
rect 24668 31668 24724 31726
rect 24668 30548 24724 31612
rect 25340 31668 25396 31678
rect 25340 31574 25396 31612
rect 25004 31556 25060 31566
rect 25004 31462 25060 31500
rect 24668 30482 24724 30492
rect 24556 30258 24612 30268
rect 25116 29540 25172 29550
rect 24220 28754 24500 28756
rect 24220 28702 24222 28754
rect 24274 28702 24500 28754
rect 24220 28700 24500 28702
rect 24668 28756 24724 28766
rect 24220 28690 24276 28700
rect 24108 28418 24164 28430
rect 24108 28366 24110 28418
rect 24162 28366 24164 28418
rect 24108 28308 24164 28366
rect 24108 28242 24164 28252
rect 24332 28418 24388 28430
rect 24332 28366 24334 28418
rect 24386 28366 24388 28418
rect 23772 27346 23828 27356
rect 24332 27412 24388 28366
rect 24332 27346 24388 27356
rect 24668 27188 24724 28700
rect 24892 28642 24948 28654
rect 24892 28590 24894 28642
rect 24946 28590 24948 28642
rect 24780 28420 24836 28430
rect 24892 28420 24948 28590
rect 24836 28364 24948 28420
rect 24780 28354 24836 28364
rect 24220 27186 24724 27188
rect 24220 27134 24670 27186
rect 24722 27134 24724 27186
rect 24220 27132 24724 27134
rect 24108 27076 24164 27086
rect 23996 26068 24052 26078
rect 23884 26066 24052 26068
rect 23884 26014 23998 26066
rect 24050 26014 24052 26066
rect 23884 26012 24052 26014
rect 23884 25618 23940 26012
rect 23996 26002 24052 26012
rect 23884 25566 23886 25618
rect 23938 25566 23940 25618
rect 23884 25508 23940 25566
rect 23884 25442 23940 25452
rect 23772 25396 23828 25406
rect 23772 25302 23828 25340
rect 23660 24892 23828 24948
rect 23772 24052 23828 24892
rect 23772 23986 23828 23996
rect 23884 24164 23940 24174
rect 24108 24164 24164 27020
rect 24220 27074 24276 27132
rect 24668 27122 24724 27132
rect 24220 27022 24222 27074
rect 24274 27022 24276 27074
rect 24220 27010 24276 27022
rect 24332 26628 24388 26638
rect 24332 26290 24388 26572
rect 24332 26238 24334 26290
rect 24386 26238 24388 26290
rect 24332 26226 24388 26238
rect 24556 26180 24612 26190
rect 24444 26178 24612 26180
rect 24444 26126 24558 26178
rect 24610 26126 24612 26178
rect 24444 26124 24612 26126
rect 24332 25732 24388 25742
rect 24444 25732 24500 26124
rect 24556 26114 24612 26124
rect 24332 25730 24500 25732
rect 24332 25678 24334 25730
rect 24386 25678 24500 25730
rect 24332 25676 24500 25678
rect 24332 25666 24388 25676
rect 24780 25508 24836 25518
rect 24780 25414 24836 25452
rect 24220 25396 24276 25406
rect 24220 25302 24276 25340
rect 25004 25282 25060 25294
rect 25004 25230 25006 25282
rect 25058 25230 25060 25282
rect 25004 24724 25060 25230
rect 25004 24658 25060 24668
rect 23884 24162 24164 24164
rect 23884 24110 23886 24162
rect 23938 24110 24164 24162
rect 23884 24108 24164 24110
rect 22988 22430 22990 22482
rect 23042 22430 23044 22482
rect 22988 22418 23044 22430
rect 23212 23266 23380 23268
rect 23212 23214 23326 23266
rect 23378 23214 23380 23266
rect 23212 23212 23380 23214
rect 22092 21858 22148 21868
rect 23100 21924 23156 21934
rect 22988 21476 23044 21486
rect 21532 20974 21534 21026
rect 21586 20974 21588 21026
rect 21532 20962 21588 20974
rect 21644 21196 21812 21252
rect 21868 21474 23044 21476
rect 21868 21422 22990 21474
rect 23042 21422 23044 21474
rect 21868 21420 23044 21422
rect 21644 20244 21700 21196
rect 21868 21026 21924 21420
rect 22988 21410 23044 21420
rect 21868 20974 21870 21026
rect 21922 20974 21924 21026
rect 21868 20962 21924 20974
rect 21756 20804 21812 20814
rect 21756 20710 21812 20748
rect 21420 20076 21588 20132
rect 21196 19966 21198 20018
rect 21250 19966 21252 20018
rect 21196 19954 21252 19966
rect 20748 19740 21140 19796
rect 21420 19906 21476 19918
rect 21420 19854 21422 19906
rect 21474 19854 21476 19906
rect 20748 19458 20804 19740
rect 20748 19406 20750 19458
rect 20802 19406 20804 19458
rect 20748 19394 20804 19406
rect 20524 18386 20580 18396
rect 19516 17726 19518 17778
rect 19570 17726 19572 17778
rect 19516 17714 19572 17726
rect 19628 17892 19684 17902
rect 19628 17668 19684 17836
rect 19740 17668 19796 17678
rect 19628 17666 19796 17668
rect 19628 17614 19742 17666
rect 19794 17614 19796 17666
rect 19628 17612 19796 17614
rect 19516 17556 19572 17566
rect 19404 17554 19572 17556
rect 19404 17502 19518 17554
rect 19570 17502 19572 17554
rect 19404 17500 19572 17502
rect 19516 17490 19572 17500
rect 19628 16882 19684 17612
rect 19740 17602 19796 17612
rect 20076 17666 20132 17678
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 20076 17444 20132 17614
rect 20076 17388 20244 17444
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 17108 20244 17388
rect 19628 16830 19630 16882
rect 19682 16830 19684 16882
rect 19628 16818 19684 16830
rect 20076 17052 20244 17108
rect 19292 16770 19572 16772
rect 19292 16718 19294 16770
rect 19346 16718 19572 16770
rect 19292 16716 19572 16718
rect 19292 16706 19348 16716
rect 18844 16660 18900 16670
rect 18844 16658 19012 16660
rect 18844 16606 18846 16658
rect 18898 16606 19012 16658
rect 18844 16604 19012 16606
rect 18844 16594 18900 16604
rect 18564 14924 18676 14980
rect 18732 16212 18788 16222
rect 18732 15090 18788 16156
rect 18956 16098 19012 16604
rect 18956 16046 18958 16098
rect 19010 16046 19012 16098
rect 18956 16034 19012 16046
rect 19516 16100 19572 16716
rect 19292 15876 19348 15886
rect 19292 15782 19348 15820
rect 19068 15316 19124 15326
rect 19068 15222 19124 15260
rect 19404 15314 19460 15326
rect 19404 15262 19406 15314
rect 19458 15262 19460 15314
rect 18732 15038 18734 15090
rect 18786 15038 18788 15090
rect 18508 14914 18564 14924
rect 18396 14868 18452 14878
rect 18396 14530 18452 14812
rect 18732 14754 18788 15038
rect 18956 15202 19012 15214
rect 18956 15150 18958 15202
rect 19010 15150 19012 15202
rect 18956 14980 19012 15150
rect 18956 14914 19012 14924
rect 18732 14702 18734 14754
rect 18786 14702 18788 14754
rect 18732 14690 18788 14702
rect 18956 14756 19012 14766
rect 18396 14478 18398 14530
rect 18450 14478 18452 14530
rect 18396 14308 18452 14478
rect 18956 14530 19012 14700
rect 19292 14532 19348 14542
rect 18956 14478 18958 14530
rect 19010 14478 19012 14530
rect 18956 14466 19012 14478
rect 19068 14530 19348 14532
rect 19068 14478 19294 14530
rect 19346 14478 19348 14530
rect 19068 14476 19348 14478
rect 18396 14242 18452 14252
rect 18620 14306 18676 14318
rect 19068 14308 19124 14476
rect 19292 14420 19348 14476
rect 19292 14354 19348 14364
rect 18620 14254 18622 14306
rect 18674 14254 18676 14306
rect 18284 13878 18340 13916
rect 18172 13806 18174 13858
rect 18226 13806 18228 13858
rect 18172 13524 18228 13806
rect 18172 13458 18228 13468
rect 17948 13300 18004 13310
rect 17836 12180 17892 12190
rect 17836 12086 17892 12124
rect 17948 12178 18004 13244
rect 17948 12126 17950 12178
rect 18002 12126 18004 12178
rect 17836 11844 17892 11854
rect 17724 11788 17836 11844
rect 17836 11778 17892 11788
rect 17612 11620 17668 11630
rect 17948 11620 18004 12126
rect 17612 11526 17668 11564
rect 17724 11564 18004 11620
rect 17612 11396 17668 11406
rect 17724 11396 17780 11564
rect 17612 11394 17780 11396
rect 17612 11342 17614 11394
rect 17666 11342 17780 11394
rect 17612 11340 17780 11342
rect 17836 11396 17892 11406
rect 17612 11330 17668 11340
rect 17836 11302 17892 11340
rect 17948 11284 18004 11294
rect 18060 11284 18116 13356
rect 18508 12068 18564 12078
rect 18620 12068 18676 14254
rect 18956 14252 19124 14308
rect 19180 14306 19236 14318
rect 19180 14254 19182 14306
rect 19234 14254 19236 14306
rect 18956 13636 19012 14252
rect 19180 14196 19236 14254
rect 19180 14140 19348 14196
rect 18956 13570 19012 13580
rect 19068 13972 19124 13982
rect 19068 13858 19124 13916
rect 19068 13806 19070 13858
rect 19122 13806 19124 13858
rect 18732 12962 18788 12974
rect 18732 12910 18734 12962
rect 18786 12910 18788 12962
rect 18732 12404 18788 12910
rect 19068 12962 19124 13806
rect 19180 13860 19236 13870
rect 19180 13766 19236 13804
rect 19292 13748 19348 14140
rect 19404 13970 19460 15262
rect 19404 13918 19406 13970
rect 19458 13918 19460 13970
rect 19404 13906 19460 13918
rect 19516 13748 19572 16044
rect 20076 15988 20132 17052
rect 20076 15876 20132 15932
rect 20076 15820 20244 15876
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19740 15540 19796 15550
rect 20188 15540 20244 15820
rect 19740 15446 19796 15484
rect 20076 15484 20244 15540
rect 19628 15316 19684 15354
rect 19628 15250 19684 15260
rect 19852 15314 19908 15326
rect 19852 15262 19854 15314
rect 19906 15262 19908 15314
rect 19740 14420 19796 14430
rect 19852 14420 19908 15262
rect 19796 14364 19908 14420
rect 19964 15314 20020 15326
rect 19964 15262 19966 15314
rect 20018 15262 20020 15314
rect 19964 14980 20020 15262
rect 19740 14326 19796 14364
rect 19964 14308 20020 14924
rect 20076 14530 20132 15484
rect 20860 15148 20916 19740
rect 21420 19458 21476 19854
rect 21420 19406 21422 19458
rect 21474 19406 21476 19458
rect 21420 19394 21476 19406
rect 21532 19124 21588 20076
rect 21644 20130 21700 20188
rect 21644 20078 21646 20130
rect 21698 20078 21700 20130
rect 21644 19460 21700 20078
rect 21756 20132 21812 20142
rect 21756 20020 21812 20076
rect 21868 20020 21924 20030
rect 21756 20018 21924 20020
rect 21756 19966 21870 20018
rect 21922 19966 21924 20018
rect 21756 19964 21924 19966
rect 21868 19954 21924 19964
rect 21644 19394 21700 19404
rect 21756 19346 21812 19358
rect 21756 19294 21758 19346
rect 21810 19294 21812 19346
rect 21644 19124 21700 19134
rect 21308 19122 21700 19124
rect 21308 19070 21646 19122
rect 21698 19070 21700 19122
rect 21308 19068 21700 19070
rect 20972 18676 21028 18686
rect 20972 18582 21028 18620
rect 20860 15092 21140 15148
rect 20076 14478 20078 14530
rect 20130 14478 20132 14530
rect 20076 14466 20132 14478
rect 20748 14868 20804 14878
rect 20748 14530 20804 14812
rect 20748 14478 20750 14530
rect 20802 14478 20804 14530
rect 20412 14308 20468 14318
rect 19964 14306 20468 14308
rect 19964 14254 20414 14306
rect 20466 14254 20468 14306
rect 19964 14252 20468 14254
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20300 14084 20356 14094
rect 20300 13970 20356 14028
rect 20300 13918 20302 13970
rect 20354 13918 20356 13970
rect 20300 13906 20356 13918
rect 19852 13748 19908 13758
rect 19292 13746 19908 13748
rect 19292 13694 19854 13746
rect 19906 13694 19908 13746
rect 19292 13692 19908 13694
rect 19852 13682 19908 13692
rect 19516 13524 19572 13534
rect 19516 12964 19572 13468
rect 20412 13412 20468 14252
rect 20748 14196 20804 14478
rect 20748 14130 20804 14140
rect 20748 13972 20804 13982
rect 20748 13878 20804 13916
rect 19068 12910 19070 12962
rect 19122 12910 19124 12962
rect 19068 12898 19124 12910
rect 19180 12962 19572 12964
rect 19180 12910 19518 12962
rect 19570 12910 19572 12962
rect 19180 12908 19572 12910
rect 18956 12404 19012 12414
rect 18732 12348 18956 12404
rect 18956 12310 19012 12348
rect 19180 12180 19236 12908
rect 19516 12898 19572 12908
rect 20300 13356 20468 13412
rect 18564 12012 18676 12068
rect 18956 12124 19236 12180
rect 19292 12738 19348 12750
rect 19292 12686 19294 12738
rect 19346 12686 19348 12738
rect 18508 12002 18564 12012
rect 18732 11844 18788 11854
rect 18172 11732 18228 11742
rect 18172 11508 18228 11676
rect 18620 11508 18676 11518
rect 18172 11506 18676 11508
rect 18172 11454 18622 11506
rect 18674 11454 18676 11506
rect 18172 11452 18676 11454
rect 18172 11394 18228 11452
rect 18620 11442 18676 11452
rect 18172 11342 18174 11394
rect 18226 11342 18228 11394
rect 18172 11330 18228 11342
rect 18004 11228 18116 11284
rect 17948 11218 18004 11228
rect 16044 9886 16046 9938
rect 16098 9886 16100 9938
rect 16044 9874 16100 9886
rect 17052 10220 17556 10276
rect 15372 9826 15428 9838
rect 15372 9774 15374 9826
rect 15426 9774 15428 9826
rect 14700 8878 14702 8930
rect 14754 8878 14756 8930
rect 14700 8148 14756 8878
rect 14700 8082 14756 8092
rect 14924 9042 14980 9054
rect 14924 8990 14926 9042
rect 14978 8990 14980 9042
rect 14364 7982 14366 8034
rect 14418 7982 14420 8034
rect 14364 7812 14420 7982
rect 14364 7746 14420 7756
rect 14924 7700 14980 8990
rect 15372 8484 15428 9774
rect 15372 8418 15428 8428
rect 16380 8484 16436 8494
rect 16380 8258 16436 8428
rect 17052 8370 17108 10220
rect 18172 9938 18228 9950
rect 18172 9886 18174 9938
rect 18226 9886 18228 9938
rect 18172 9716 18228 9886
rect 18620 9940 18676 9950
rect 18732 9940 18788 11788
rect 18956 11282 19012 12124
rect 19292 12068 19348 12686
rect 19404 12738 19460 12750
rect 19404 12686 19406 12738
rect 19458 12686 19460 12738
rect 19404 12180 19460 12686
rect 19628 12738 19684 12750
rect 19628 12686 19630 12738
rect 19682 12686 19684 12738
rect 19404 12114 19460 12124
rect 19516 12628 19572 12638
rect 19292 12002 19348 12012
rect 19516 11620 19572 12572
rect 19628 12292 19684 12686
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19740 12292 19796 12302
rect 19628 12236 19740 12292
rect 19740 12226 19796 12236
rect 20300 12292 20356 13356
rect 21084 13188 21140 15092
rect 21308 13412 21364 19068
rect 21644 19058 21700 19068
rect 21532 18450 21588 18462
rect 21532 18398 21534 18450
rect 21586 18398 21588 18450
rect 21532 17780 21588 18398
rect 21756 18452 21812 19294
rect 22204 18452 22260 18462
rect 21756 18450 22260 18452
rect 21756 18398 22206 18450
rect 22258 18398 22260 18450
rect 21756 18396 22260 18398
rect 22204 18386 22260 18396
rect 21532 16884 21588 17724
rect 21532 16828 21924 16884
rect 21868 15314 21924 16828
rect 22316 16212 22372 16222
rect 22092 15986 22148 15998
rect 22092 15934 22094 15986
rect 22146 15934 22148 15986
rect 22092 15540 22148 15934
rect 22316 15986 22372 16156
rect 22316 15934 22318 15986
rect 22370 15934 22372 15986
rect 22316 15922 22372 15934
rect 22428 16210 22484 16222
rect 22428 16158 22430 16210
rect 22482 16158 22484 16210
rect 22092 15474 22148 15484
rect 22428 15428 22484 16158
rect 22876 16212 22932 16222
rect 22876 16118 22932 16156
rect 23100 15652 23156 21868
rect 23100 15586 23156 15596
rect 23212 17444 23268 23212
rect 23324 23202 23380 23212
rect 23660 23938 23716 23950
rect 23660 23886 23662 23938
rect 23714 23886 23716 23938
rect 23660 19236 23716 23886
rect 23772 21586 23828 21598
rect 23772 21534 23774 21586
rect 23826 21534 23828 21586
rect 23772 21476 23828 21534
rect 23772 21410 23828 21420
rect 23884 20804 23940 24108
rect 24220 23940 24276 23950
rect 24220 23846 24276 23884
rect 24444 23826 24500 23838
rect 24444 23774 24446 23826
rect 24498 23774 24500 23826
rect 24332 23714 24388 23726
rect 24332 23662 24334 23714
rect 24386 23662 24388 23714
rect 24332 22708 24388 23662
rect 24444 23268 24500 23774
rect 24444 23202 24500 23212
rect 25116 23156 25172 29484
rect 25228 28756 25284 28766
rect 25228 28642 25284 28700
rect 25228 28590 25230 28642
rect 25282 28590 25284 28642
rect 25228 28578 25284 28590
rect 25452 28308 25508 34076
rect 25788 33234 25844 33246
rect 25788 33182 25790 33234
rect 25842 33182 25844 33234
rect 25676 32788 25732 32798
rect 25788 32788 25844 33182
rect 25676 32786 25844 32788
rect 25676 32734 25678 32786
rect 25730 32734 25844 32786
rect 25676 32732 25844 32734
rect 25676 32722 25732 32732
rect 25564 32562 25620 32574
rect 25564 32510 25566 32562
rect 25618 32510 25620 32562
rect 25564 32452 25620 32510
rect 25788 32564 25844 32574
rect 25788 32470 25844 32508
rect 25900 32452 25956 34188
rect 26012 32788 26068 34412
rect 26124 34130 26180 34142
rect 26124 34078 26126 34130
rect 26178 34078 26180 34130
rect 26124 32788 26180 34078
rect 26236 34132 26292 34862
rect 26572 34916 26628 35084
rect 26684 34916 26740 34926
rect 26572 34914 26740 34916
rect 26572 34862 26686 34914
rect 26738 34862 26740 34914
rect 26572 34860 26740 34862
rect 26684 34850 26740 34860
rect 26236 34066 26292 34076
rect 26124 32732 26292 32788
rect 26012 32676 26068 32732
rect 26012 32620 26180 32676
rect 26012 32452 26068 32462
rect 25900 32396 26012 32452
rect 25564 32386 25620 32396
rect 26012 32386 26068 32396
rect 25900 31556 25956 31566
rect 25788 31554 25956 31556
rect 25788 31502 25902 31554
rect 25954 31502 25956 31554
rect 25788 31500 25956 31502
rect 25452 28242 25508 28252
rect 25564 30994 25620 31006
rect 25564 30942 25566 30994
rect 25618 30942 25620 30994
rect 25340 27746 25396 27758
rect 25340 27694 25342 27746
rect 25394 27694 25396 27746
rect 25340 27412 25396 27694
rect 25340 27346 25396 27356
rect 25564 24836 25620 30942
rect 25676 30996 25732 31006
rect 25788 30996 25844 31500
rect 25900 31490 25956 31500
rect 25732 30940 25844 30996
rect 25900 31106 25956 31118
rect 25900 31054 25902 31106
rect 25954 31054 25956 31106
rect 25676 30930 25732 30940
rect 25900 30884 25956 31054
rect 25788 30828 25956 30884
rect 25788 30212 25844 30828
rect 26012 30772 26068 30782
rect 25788 30146 25844 30156
rect 25900 30716 26012 30772
rect 25900 30210 25956 30716
rect 26012 30706 26068 30716
rect 25900 30158 25902 30210
rect 25954 30158 25956 30210
rect 25900 30146 25956 30158
rect 26012 29988 26068 29998
rect 25900 29986 26068 29988
rect 25900 29934 26014 29986
rect 26066 29934 26068 29986
rect 25900 29932 26068 29934
rect 25900 28754 25956 29932
rect 26012 29922 26068 29932
rect 25900 28702 25902 28754
rect 25954 28702 25956 28754
rect 25900 28690 25956 28702
rect 25788 28308 25844 28318
rect 25788 27186 25844 28252
rect 25788 27134 25790 27186
rect 25842 27134 25844 27186
rect 25788 27122 25844 27134
rect 25564 24770 25620 24780
rect 25788 24724 25844 24734
rect 25788 24630 25844 24668
rect 26124 24722 26180 32620
rect 26236 31780 26292 32732
rect 26908 32786 26964 35532
rect 27244 35026 27300 36204
rect 28476 36260 28532 36270
rect 27244 34974 27246 35026
rect 27298 34974 27300 35026
rect 27244 34962 27300 34974
rect 27692 35252 27748 35262
rect 26908 32734 26910 32786
rect 26962 32734 26964 32786
rect 26236 31332 26292 31724
rect 26572 31780 26628 31790
rect 26572 31686 26628 31724
rect 26236 31266 26292 31276
rect 26684 31554 26740 31566
rect 26684 31502 26686 31554
rect 26738 31502 26740 31554
rect 26460 31220 26516 31230
rect 26684 31220 26740 31502
rect 26796 31556 26852 31566
rect 26796 31462 26852 31500
rect 26460 31218 26740 31220
rect 26460 31166 26462 31218
rect 26514 31166 26740 31218
rect 26460 31164 26740 31166
rect 26908 31218 26964 32734
rect 27356 32788 27412 32798
rect 27356 32694 27412 32732
rect 26908 31166 26910 31218
rect 26962 31166 26964 31218
rect 26460 31154 26516 31164
rect 26908 31154 26964 31166
rect 27020 31892 27076 31902
rect 26236 31108 26292 31118
rect 26236 31014 26292 31052
rect 26796 30994 26852 31006
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26572 30772 26628 30810
rect 26572 30706 26628 30716
rect 26572 30548 26628 30558
rect 26460 30212 26516 30222
rect 26460 30118 26516 30156
rect 26236 30100 26292 30110
rect 26236 30098 26404 30100
rect 26236 30046 26238 30098
rect 26290 30046 26404 30098
rect 26236 30044 26404 30046
rect 26236 30034 26292 30044
rect 26348 29204 26404 30044
rect 26572 29538 26628 30492
rect 26796 30212 26852 30942
rect 26796 30146 26852 30156
rect 26908 30100 26964 30110
rect 26908 30006 26964 30044
rect 27020 29764 27076 31836
rect 27580 31892 27636 31902
rect 27132 31778 27188 31790
rect 27132 31726 27134 31778
rect 27186 31726 27188 31778
rect 27132 31668 27188 31726
rect 27580 31778 27636 31836
rect 27580 31726 27582 31778
rect 27634 31726 27636 31778
rect 27580 31714 27636 31726
rect 27468 31668 27524 31678
rect 27132 31666 27524 31668
rect 27132 31614 27470 31666
rect 27522 31614 27524 31666
rect 27132 31612 27524 31614
rect 27244 31218 27300 31230
rect 27244 31166 27246 31218
rect 27298 31166 27300 31218
rect 27244 30994 27300 31166
rect 27244 30942 27246 30994
rect 27298 30942 27300 30994
rect 27132 30212 27188 30222
rect 27132 30118 27188 30156
rect 26572 29486 26574 29538
rect 26626 29486 26628 29538
rect 26572 29428 26628 29486
rect 26908 29708 27076 29764
rect 27132 29988 27188 29998
rect 26908 29538 26964 29708
rect 26908 29486 26910 29538
rect 26962 29486 26964 29538
rect 26572 29362 26628 29372
rect 26684 29426 26740 29438
rect 26684 29374 26686 29426
rect 26738 29374 26740 29426
rect 26684 29204 26740 29374
rect 26348 29148 26740 29204
rect 26908 28532 26964 29486
rect 27020 29540 27076 29550
rect 27132 29540 27188 29932
rect 27076 29484 27188 29540
rect 27020 29446 27076 29484
rect 26908 28466 26964 28476
rect 27244 27860 27300 30942
rect 27468 30436 27524 31612
rect 27580 30436 27636 30446
rect 27468 30434 27636 30436
rect 27468 30382 27582 30434
rect 27634 30382 27636 30434
rect 27468 30380 27636 30382
rect 27580 30370 27636 30380
rect 27692 30212 27748 35196
rect 27916 33458 27972 33470
rect 27916 33406 27918 33458
rect 27970 33406 27972 33458
rect 27916 33236 27972 33406
rect 28476 33460 28532 36204
rect 28588 34692 28644 37884
rect 29148 37828 29204 39342
rect 29372 38162 29428 39564
rect 29820 39396 29876 39406
rect 29820 39058 29876 39340
rect 29820 39006 29822 39058
rect 29874 39006 29876 39058
rect 29820 38994 29876 39006
rect 29932 39394 29988 39406
rect 29932 39342 29934 39394
rect 29986 39342 29988 39394
rect 29932 38724 29988 39342
rect 30044 39394 30100 39406
rect 30044 39342 30046 39394
rect 30098 39342 30100 39394
rect 30044 38834 30100 39342
rect 30044 38782 30046 38834
rect 30098 38782 30100 38834
rect 30044 38770 30100 38782
rect 30156 39394 30212 39406
rect 30156 39342 30158 39394
rect 30210 39342 30212 39394
rect 30156 38836 30212 39342
rect 29932 38658 29988 38668
rect 29372 38110 29374 38162
rect 29426 38110 29428 38162
rect 29372 38098 29428 38110
rect 30156 38164 30212 38780
rect 30156 38070 30212 38108
rect 30268 38612 30324 40908
rect 30380 40898 30436 40908
rect 30828 40962 30884 40974
rect 30828 40910 30830 40962
rect 30882 40910 30884 40962
rect 30380 40292 30436 40302
rect 30380 40198 30436 40236
rect 30828 39618 30884 40910
rect 40124 40964 40180 40974
rect 40124 40962 40292 40964
rect 40124 40910 40126 40962
rect 40178 40910 40292 40962
rect 40124 40908 40292 40910
rect 40124 40898 40180 40908
rect 40124 40514 40180 40526
rect 40124 40462 40126 40514
rect 40178 40462 40180 40514
rect 31948 40292 32004 40302
rect 31164 39732 31220 39742
rect 31836 39732 31892 39742
rect 31164 39730 31892 39732
rect 31164 39678 31166 39730
rect 31218 39678 31838 39730
rect 31890 39678 31892 39730
rect 31164 39676 31892 39678
rect 31164 39666 31220 39676
rect 31836 39666 31892 39676
rect 31948 39730 32004 40236
rect 32508 40292 32564 40302
rect 32508 40290 32788 40292
rect 32508 40238 32510 40290
rect 32562 40238 32788 40290
rect 32508 40236 32788 40238
rect 32508 40226 32564 40236
rect 31948 39678 31950 39730
rect 32002 39678 32004 39730
rect 31948 39666 32004 39678
rect 30828 39566 30830 39618
rect 30882 39566 30884 39618
rect 29148 37268 29204 37772
rect 29148 37202 29204 37212
rect 29708 38050 29764 38062
rect 29708 37998 29710 38050
rect 29762 37998 29764 38050
rect 29708 37940 29764 37998
rect 29148 36596 29204 36606
rect 29148 36370 29204 36540
rect 29708 36596 29764 37884
rect 30268 37828 30324 38556
rect 30268 37762 30324 37772
rect 30380 39394 30436 39406
rect 30380 39342 30382 39394
rect 30434 39342 30436 39394
rect 30380 37716 30436 39342
rect 30828 38052 30884 39566
rect 32732 39620 32788 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 40124 39732 40180 40462
rect 40236 40404 40292 40908
rect 40348 40404 40404 40414
rect 40236 40348 40348 40404
rect 40348 40338 40404 40348
rect 40124 39666 40180 39676
rect 32732 39618 33124 39620
rect 32732 39566 32734 39618
rect 32786 39566 33124 39618
rect 32732 39564 33124 39566
rect 32732 39554 32788 39564
rect 31500 39506 31556 39518
rect 31500 39454 31502 39506
rect 31554 39454 31556 39506
rect 31052 39394 31108 39406
rect 31052 39342 31054 39394
rect 31106 39342 31108 39394
rect 31052 39172 31108 39342
rect 31276 39396 31332 39406
rect 31276 39302 31332 39340
rect 30940 39116 31108 39172
rect 30940 38948 30996 39116
rect 30940 38834 30996 38892
rect 30940 38782 30942 38834
rect 30994 38782 30996 38834
rect 30940 38770 30996 38782
rect 31388 38946 31444 38958
rect 31388 38894 31390 38946
rect 31442 38894 31444 38946
rect 31052 38164 31108 38174
rect 31052 38052 31108 38108
rect 31164 38052 31220 38062
rect 31052 38050 31220 38052
rect 31052 37998 31166 38050
rect 31218 37998 31220 38050
rect 31052 37996 31220 37998
rect 30828 37986 30884 37996
rect 31164 37986 31220 37996
rect 30492 37940 30548 37950
rect 30492 37846 30548 37884
rect 30940 37940 30996 37950
rect 30940 37938 31108 37940
rect 30940 37886 30942 37938
rect 30994 37886 31108 37938
rect 30940 37884 31108 37886
rect 30940 37874 30996 37884
rect 30604 37828 30660 37838
rect 30660 37772 30772 37828
rect 30604 37734 30660 37772
rect 30380 37660 30548 37716
rect 30492 37492 30548 37660
rect 30604 37492 30660 37502
rect 30492 37490 30660 37492
rect 30492 37438 30606 37490
rect 30658 37438 30660 37490
rect 30492 37436 30660 37438
rect 30604 37426 30660 37436
rect 30380 37380 30436 37390
rect 30380 37286 30436 37324
rect 30268 37268 30324 37278
rect 30268 37174 30324 37212
rect 30716 37266 30772 37772
rect 31052 37492 31108 37884
rect 31276 37492 31332 37502
rect 31052 37490 31332 37492
rect 31052 37438 31278 37490
rect 31330 37438 31332 37490
rect 31052 37436 31332 37438
rect 31388 37492 31444 38894
rect 31500 38668 31556 39454
rect 32060 39508 32116 39518
rect 32060 39414 32116 39452
rect 32508 39394 32564 39406
rect 32508 39342 32510 39394
rect 32562 39342 32564 39394
rect 32060 38948 32116 38958
rect 32060 38854 32116 38892
rect 32396 38836 32452 38846
rect 32508 38836 32564 39342
rect 32396 38834 32564 38836
rect 32396 38782 32398 38834
rect 32450 38782 32564 38834
rect 32396 38780 32564 38782
rect 32732 38948 32788 38958
rect 31724 38724 31780 38734
rect 31500 38612 31668 38668
rect 31612 38546 31668 38556
rect 31500 38500 31556 38510
rect 31500 38274 31556 38444
rect 31500 38222 31502 38274
rect 31554 38222 31556 38274
rect 31500 38210 31556 38222
rect 31724 38274 31780 38668
rect 31724 38222 31726 38274
rect 31778 38222 31780 38274
rect 31724 38210 31780 38222
rect 31836 37826 31892 37838
rect 31836 37774 31838 37826
rect 31890 37774 31892 37826
rect 31388 37436 31556 37492
rect 31276 37426 31332 37436
rect 31500 37380 31556 37436
rect 31500 37314 31556 37324
rect 30716 37214 30718 37266
rect 30770 37214 30772 37266
rect 30716 37202 30772 37214
rect 31052 37268 31108 37278
rect 31164 37268 31220 37278
rect 31108 37266 31220 37268
rect 31108 37214 31166 37266
rect 31218 37214 31220 37266
rect 31108 37212 31220 37214
rect 29708 36530 29764 36540
rect 29148 36318 29150 36370
rect 29202 36318 29204 36370
rect 29148 36306 29204 36318
rect 29372 36482 29428 36494
rect 29372 36430 29374 36482
rect 29426 36430 29428 36482
rect 28588 34626 28644 34636
rect 29036 34132 29092 34142
rect 29260 34132 29316 34142
rect 29036 34130 29260 34132
rect 29036 34078 29038 34130
rect 29090 34078 29260 34130
rect 29036 34076 29260 34078
rect 29036 34066 29092 34076
rect 28476 33366 28532 33404
rect 27916 33170 27972 33180
rect 28924 33012 28980 33022
rect 28140 32788 28196 32798
rect 27804 31892 27860 31902
rect 27804 30434 27860 31836
rect 28140 31778 28196 32732
rect 28924 32674 28980 32956
rect 28924 32622 28926 32674
rect 28978 32622 28980 32674
rect 28924 32610 28980 32622
rect 29036 32564 29092 32574
rect 29036 32470 29092 32508
rect 28140 31726 28142 31778
rect 28194 31726 28196 31778
rect 28140 31714 28196 31726
rect 27804 30382 27806 30434
rect 27858 30382 27860 30434
rect 27804 30370 27860 30382
rect 28028 31556 28084 31566
rect 27468 30156 27748 30212
rect 28028 30210 28084 31500
rect 28028 30158 28030 30210
rect 28082 30158 28084 30210
rect 27356 27972 27412 27982
rect 27356 27878 27412 27916
rect 27244 27794 27300 27804
rect 27244 27636 27300 27646
rect 26684 27634 27300 27636
rect 26684 27582 27246 27634
rect 27298 27582 27300 27634
rect 26684 27580 27300 27582
rect 27468 27636 27524 30156
rect 28028 30146 28084 30158
rect 28364 30548 28420 30558
rect 28364 30210 28420 30492
rect 28364 30158 28366 30210
rect 28418 30158 28420 30210
rect 28364 30146 28420 30158
rect 28252 30100 28308 30110
rect 28028 28754 28084 28766
rect 28028 28702 28030 28754
rect 28082 28702 28084 28754
rect 27916 28532 27972 28542
rect 27916 27970 27972 28476
rect 27916 27918 27918 27970
rect 27970 27918 27972 27970
rect 27580 27858 27636 27870
rect 27580 27806 27582 27858
rect 27634 27806 27636 27858
rect 27580 27748 27636 27806
rect 27916 27860 27972 27918
rect 28028 27860 28084 28702
rect 28252 28532 28308 30044
rect 28476 29986 28532 29998
rect 28476 29934 28478 29986
rect 28530 29934 28532 29986
rect 28476 29652 28532 29934
rect 28700 29988 28756 29998
rect 29148 29988 29204 34076
rect 29260 34066 29316 34076
rect 29372 34130 29428 36430
rect 30380 36260 30436 36270
rect 30380 35810 30436 36204
rect 30380 35758 30382 35810
rect 30434 35758 30436 35810
rect 30380 35746 30436 35758
rect 30940 35476 30996 35486
rect 30828 35474 30996 35476
rect 30828 35422 30942 35474
rect 30994 35422 30996 35474
rect 30828 35420 30996 35422
rect 30828 34914 30884 35420
rect 30940 35410 30996 35420
rect 31052 35140 31108 37212
rect 31164 37202 31220 37212
rect 31388 37266 31444 37278
rect 31388 37214 31390 37266
rect 31442 37214 31444 37266
rect 31388 37044 31444 37214
rect 31388 36978 31444 36988
rect 31724 37268 31780 37278
rect 31276 36260 31332 36270
rect 31332 36204 31668 36260
rect 31276 36166 31332 36204
rect 31500 35812 31556 35822
rect 31500 35718 31556 35756
rect 31276 35700 31332 35710
rect 31276 35606 31332 35644
rect 31052 35074 31108 35084
rect 31164 35476 31220 35486
rect 30828 34862 30830 34914
rect 30882 34862 30884 34914
rect 30828 34850 30884 34862
rect 30492 34804 30548 34814
rect 30492 34710 30548 34748
rect 31164 34804 31220 35420
rect 31612 34914 31668 36204
rect 31612 34862 31614 34914
rect 31666 34862 31668 34914
rect 31612 34850 31668 34862
rect 29932 34692 29988 34702
rect 29372 34078 29374 34130
rect 29426 34078 29428 34130
rect 29260 33234 29316 33246
rect 29260 33182 29262 33234
rect 29314 33182 29316 33234
rect 29260 32564 29316 33182
rect 29260 32470 29316 32508
rect 29372 31668 29428 34078
rect 29708 34242 29764 34254
rect 29708 34190 29710 34242
rect 29762 34190 29764 34242
rect 29708 33348 29764 34190
rect 29708 33282 29764 33292
rect 29932 33236 29988 34636
rect 30156 34690 30212 34702
rect 30156 34638 30158 34690
rect 30210 34638 30212 34690
rect 30156 34580 30212 34638
rect 30156 34514 30212 34524
rect 30380 34690 30436 34702
rect 30380 34638 30382 34690
rect 30434 34638 30436 34690
rect 30268 34242 30324 34254
rect 30268 34190 30270 34242
rect 30322 34190 30324 34242
rect 30156 34132 30212 34142
rect 30156 34038 30212 34076
rect 30268 33684 30324 34190
rect 30156 33628 30324 33684
rect 30156 33460 30212 33628
rect 30380 33572 30436 34638
rect 31052 34692 31108 34702
rect 31164 34692 31220 34748
rect 31052 34690 31220 34692
rect 31052 34638 31054 34690
rect 31106 34638 31220 34690
rect 31052 34636 31220 34638
rect 31052 34626 31108 34636
rect 30492 34356 30548 34394
rect 30492 34290 30548 34300
rect 31052 34356 31108 34366
rect 31052 34242 31108 34300
rect 31052 34190 31054 34242
rect 31106 34190 31108 34242
rect 31052 34178 31108 34190
rect 30380 33506 30436 33516
rect 30492 34132 30548 34142
rect 30156 33394 30212 33404
rect 30268 33458 30324 33470
rect 30268 33406 30270 33458
rect 30322 33406 30324 33458
rect 30268 33236 30324 33406
rect 30380 33348 30436 33358
rect 30380 33254 30436 33292
rect 29932 33180 30212 33236
rect 29484 33124 29540 33134
rect 29484 32674 29540 33068
rect 29932 32788 29988 32798
rect 29484 32622 29486 32674
rect 29538 32622 29540 32674
rect 29484 32610 29540 32622
rect 29596 32786 29988 32788
rect 29596 32734 29934 32786
rect 29986 32734 29988 32786
rect 29596 32732 29988 32734
rect 29596 31892 29652 32732
rect 29932 32722 29988 32732
rect 29820 32562 29876 32574
rect 29820 32510 29822 32562
rect 29874 32510 29876 32562
rect 29820 31892 29876 32510
rect 30044 32562 30100 32574
rect 30044 32510 30046 32562
rect 30098 32510 30100 32562
rect 30044 32340 30100 32510
rect 30044 32274 30100 32284
rect 29820 31836 30100 31892
rect 29596 31826 29652 31836
rect 29372 31612 29764 31668
rect 29484 30548 29540 30558
rect 28700 29986 29092 29988
rect 28700 29934 28702 29986
rect 28754 29934 29092 29986
rect 28700 29932 29092 29934
rect 28700 29922 28756 29932
rect 29036 29652 29092 29932
rect 29148 29922 29204 29932
rect 29260 30210 29316 30222
rect 29260 30158 29262 30210
rect 29314 30158 29316 30210
rect 29260 29876 29316 30158
rect 29484 30098 29540 30492
rect 29484 30046 29486 30098
rect 29538 30046 29540 30098
rect 29484 30034 29540 30046
rect 29596 30100 29652 30110
rect 29260 29810 29316 29820
rect 29036 29596 29540 29652
rect 28476 29586 28532 29596
rect 29484 29538 29540 29596
rect 29596 29650 29652 30044
rect 29596 29598 29598 29650
rect 29650 29598 29652 29650
rect 29596 29586 29652 29598
rect 29484 29486 29486 29538
rect 29538 29486 29540 29538
rect 29484 29474 29540 29486
rect 29596 29204 29652 29214
rect 29484 29202 29652 29204
rect 29484 29150 29598 29202
rect 29650 29150 29652 29202
rect 29484 29148 29652 29150
rect 28476 28756 28532 28766
rect 28476 28662 28532 28700
rect 28252 28476 28532 28532
rect 28252 27860 28308 27870
rect 28028 27858 28308 27860
rect 28028 27806 28254 27858
rect 28306 27806 28308 27858
rect 28028 27804 28308 27806
rect 27916 27794 27972 27804
rect 27580 27692 27860 27748
rect 27468 27580 27748 27636
rect 26684 27186 26740 27580
rect 27244 27570 27300 27580
rect 26684 27134 26686 27186
rect 26738 27134 26740 27186
rect 26684 27122 26740 27134
rect 27692 27186 27748 27580
rect 27804 27524 27860 27692
rect 27804 27468 28084 27524
rect 27692 27134 27694 27186
rect 27746 27134 27748 27186
rect 27692 27122 27748 27134
rect 28028 27186 28084 27468
rect 28028 27134 28030 27186
rect 28082 27134 28084 27186
rect 28028 27122 28084 27134
rect 26236 27074 26292 27086
rect 26236 27022 26238 27074
rect 26290 27022 26292 27074
rect 26236 26180 26292 27022
rect 27580 27074 27636 27086
rect 27580 27022 27582 27074
rect 27634 27022 27636 27074
rect 27580 26964 27636 27022
rect 27580 26898 27636 26908
rect 27692 26292 27748 26302
rect 27692 26198 27748 26236
rect 26236 26114 26292 26124
rect 26908 26180 26964 26190
rect 26908 26086 26964 26124
rect 28252 26180 28308 27804
rect 28364 26852 28420 26862
rect 28364 26402 28420 26796
rect 28364 26350 28366 26402
rect 28418 26350 28420 26402
rect 28364 26338 28420 26350
rect 28252 26114 28308 26124
rect 26124 24670 26126 24722
rect 26178 24670 26180 24722
rect 26124 24658 26180 24670
rect 26684 24724 26740 24734
rect 26740 24668 26852 24724
rect 26684 24630 26740 24668
rect 25228 24610 25284 24622
rect 25228 24558 25230 24610
rect 25282 24558 25284 24610
rect 25228 24052 25284 24558
rect 25228 23986 25284 23996
rect 25116 23100 25284 23156
rect 24332 22652 25172 22708
rect 25116 22482 25172 22652
rect 25116 22430 25118 22482
rect 25170 22430 25172 22482
rect 25116 22418 25172 22430
rect 25228 22260 25284 23100
rect 26572 23154 26628 23166
rect 26572 23102 26574 23154
rect 26626 23102 26628 23154
rect 25116 22204 25284 22260
rect 25788 22370 25844 22382
rect 25788 22318 25790 22370
rect 25842 22318 25844 22370
rect 24220 21476 24276 21486
rect 24220 21382 24276 21420
rect 23884 20738 23940 20748
rect 24668 19572 24724 19582
rect 23772 19460 23828 19470
rect 23772 19366 23828 19404
rect 23660 19170 23716 19180
rect 24332 19236 24388 19246
rect 24332 19142 24388 19180
rect 24668 19234 24724 19516
rect 24668 19182 24670 19234
rect 24722 19182 24724 19234
rect 24668 19170 24724 19182
rect 23884 19122 23940 19134
rect 23884 19070 23886 19122
rect 23938 19070 23940 19122
rect 23884 18116 23940 19070
rect 24892 19122 24948 19134
rect 24892 19070 24894 19122
rect 24946 19070 24948 19122
rect 24780 19010 24836 19022
rect 24780 18958 24782 19010
rect 24834 18958 24836 19010
rect 24780 18452 24836 18958
rect 24780 18386 24836 18396
rect 23884 18050 23940 18060
rect 24332 18338 24388 18350
rect 24332 18286 24334 18338
rect 24386 18286 24388 18338
rect 24332 18116 24388 18286
rect 24892 18228 24948 19070
rect 25116 18340 25172 22204
rect 25340 21476 25396 21486
rect 25228 19908 25284 19918
rect 25228 19814 25284 19852
rect 24892 18162 24948 18172
rect 25004 18284 25116 18340
rect 24332 18050 24388 18060
rect 24556 17780 24612 17790
rect 24556 17686 24612 17724
rect 25004 17778 25060 18284
rect 25116 18274 25172 18284
rect 25228 19236 25284 19246
rect 25340 19236 25396 21420
rect 25788 21476 25844 22318
rect 26348 22370 26404 22382
rect 26348 22318 26350 22370
rect 26402 22318 26404 22370
rect 26348 22148 26404 22318
rect 26348 22082 26404 22092
rect 25788 21410 25844 21420
rect 26124 21476 26180 21486
rect 26124 21382 26180 21420
rect 26572 21476 26628 23102
rect 26796 22370 26852 24668
rect 27804 23492 27860 23502
rect 27860 23436 27972 23492
rect 27804 23426 27860 23436
rect 27468 23268 27524 23278
rect 27356 23042 27412 23054
rect 27356 22990 27358 23042
rect 27410 22990 27412 23042
rect 27356 22482 27412 22990
rect 27356 22430 27358 22482
rect 27410 22430 27412 22482
rect 27356 22418 27412 22430
rect 27468 22596 27524 23212
rect 26796 22318 26798 22370
rect 26850 22318 26852 22370
rect 26796 21812 26852 22318
rect 27468 22370 27524 22540
rect 27468 22318 27470 22370
rect 27522 22318 27524 22370
rect 27468 22306 27524 22318
rect 27804 23044 27860 23054
rect 27804 22370 27860 22988
rect 27804 22318 27806 22370
rect 27858 22318 27860 22370
rect 27804 22306 27860 22318
rect 26796 21746 26852 21756
rect 26908 22148 26964 22158
rect 26908 21810 26964 22092
rect 27244 22148 27300 22158
rect 27244 22054 27300 22092
rect 27916 22148 27972 23436
rect 28140 22482 28196 22494
rect 28140 22430 28142 22482
rect 28194 22430 28196 22482
rect 28028 22260 28084 22270
rect 28028 22166 28084 22204
rect 26908 21758 26910 21810
rect 26962 21758 26964 21810
rect 26908 21476 26964 21758
rect 27916 21698 27972 22092
rect 27916 21646 27918 21698
rect 27970 21646 27972 21698
rect 27916 21634 27972 21646
rect 28140 21698 28196 22430
rect 28252 22484 28308 22494
rect 28476 22484 28532 28476
rect 29036 27860 29092 27870
rect 29036 27074 29092 27804
rect 29036 27022 29038 27074
rect 29090 27022 29092 27074
rect 29036 27010 29092 27022
rect 29484 27074 29540 29148
rect 29596 29138 29652 29148
rect 29484 27022 29486 27074
rect 29538 27022 29540 27074
rect 29484 27010 29540 27022
rect 29596 27076 29652 27114
rect 29596 27010 29652 27020
rect 28588 26964 28644 27002
rect 29708 26908 29764 31612
rect 29820 31556 29876 31566
rect 29820 31462 29876 31500
rect 30044 30100 30100 31836
rect 30156 31668 30212 33180
rect 30156 31108 30212 31612
rect 30268 31332 30324 33180
rect 30492 32788 30548 34076
rect 30940 34132 30996 34142
rect 30940 34038 30996 34076
rect 31164 34020 31220 34636
rect 31276 34692 31332 34702
rect 31276 34598 31332 34636
rect 31388 34690 31444 34702
rect 31388 34638 31390 34690
rect 31442 34638 31444 34690
rect 31276 34356 31332 34366
rect 31276 34262 31332 34300
rect 31388 34242 31444 34638
rect 31388 34190 31390 34242
rect 31442 34190 31444 34242
rect 31388 34178 31444 34190
rect 30380 32732 30548 32788
rect 31052 33964 31220 34020
rect 31052 32788 31108 33964
rect 31612 33906 31668 33918
rect 31612 33854 31614 33906
rect 31666 33854 31668 33906
rect 31612 33236 31668 33854
rect 31164 33122 31220 33134
rect 31164 33070 31166 33122
rect 31218 33070 31220 33122
rect 31164 33012 31220 33070
rect 31276 33124 31332 33134
rect 31276 33030 31332 33068
rect 31388 33124 31444 33134
rect 31388 33122 31556 33124
rect 31388 33070 31390 33122
rect 31442 33070 31556 33122
rect 31388 33068 31556 33070
rect 31388 33058 31444 33068
rect 31164 32946 31220 32956
rect 31052 32732 31444 32788
rect 30380 31556 30436 32732
rect 30492 32562 30548 32574
rect 30492 32510 30494 32562
rect 30546 32510 30548 32562
rect 30492 32452 30548 32510
rect 31052 32564 31108 32574
rect 31052 32562 31332 32564
rect 31052 32510 31054 32562
rect 31106 32510 31332 32562
rect 31052 32508 31332 32510
rect 31052 32452 31108 32508
rect 30492 32396 31108 32452
rect 30828 32228 30884 32238
rect 30828 31666 30884 32172
rect 30828 31614 30830 31666
rect 30882 31614 30884 31666
rect 30828 31602 30884 31614
rect 30380 31500 30660 31556
rect 30268 31276 30548 31332
rect 30156 31042 30212 31052
rect 30044 30034 30100 30044
rect 30268 30882 30324 30894
rect 30268 30830 30270 30882
rect 30322 30830 30324 30882
rect 30268 29988 30324 30830
rect 30380 30100 30436 30110
rect 30380 30006 30436 30044
rect 30268 28756 30324 29932
rect 30380 29876 30436 29886
rect 30492 29876 30548 31276
rect 30604 30324 30660 31500
rect 30604 30258 30660 30268
rect 30716 30884 30772 30894
rect 30716 30322 30772 30828
rect 31164 30548 31220 30558
rect 30716 30270 30718 30322
rect 30770 30270 30772 30322
rect 30716 30258 30772 30270
rect 30828 30324 30884 30334
rect 30436 29820 30548 29876
rect 30604 29986 30660 29998
rect 30828 29988 30884 30268
rect 30604 29934 30606 29986
rect 30658 29934 30660 29986
rect 30380 29810 30436 29820
rect 30604 29764 30660 29934
rect 30604 29698 30660 29708
rect 30716 29986 30884 29988
rect 30716 29934 30830 29986
rect 30882 29934 30884 29986
rect 30716 29932 30884 29934
rect 30492 29652 30548 29662
rect 30492 29540 30548 29596
rect 30604 29540 30660 29550
rect 30492 29538 30660 29540
rect 30492 29486 30606 29538
rect 30658 29486 30660 29538
rect 30492 29484 30660 29486
rect 30604 29474 30660 29484
rect 30268 28690 30324 28700
rect 29820 27636 29876 27646
rect 29820 27186 29876 27580
rect 29820 27134 29822 27186
rect 29874 27134 29876 27186
rect 29820 27122 29876 27134
rect 30044 27188 30100 27198
rect 30044 27074 30100 27132
rect 30044 27022 30046 27074
rect 30098 27022 30100 27074
rect 30044 27010 30100 27022
rect 28588 26852 28756 26908
rect 28252 22370 28308 22428
rect 28252 22318 28254 22370
rect 28306 22318 28308 22370
rect 28252 22306 28308 22318
rect 28364 22428 28532 22484
rect 28588 26068 28644 26078
rect 28140 21646 28142 21698
rect 28194 21646 28196 21698
rect 27580 21588 27636 21598
rect 27580 21494 27636 21532
rect 26572 21410 26628 21420
rect 26796 21420 26964 21476
rect 27692 21474 27748 21486
rect 27692 21422 27694 21474
rect 27746 21422 27748 21474
rect 25788 20804 25844 20814
rect 25788 20242 25844 20748
rect 25788 20190 25790 20242
rect 25842 20190 25844 20242
rect 25788 20178 25844 20190
rect 26124 20132 26180 20142
rect 26124 20130 26292 20132
rect 26124 20078 26126 20130
rect 26178 20078 26292 20130
rect 26124 20076 26292 20078
rect 26124 20066 26180 20076
rect 25900 19908 25956 19918
rect 25956 19852 26180 19908
rect 25900 19842 25956 19852
rect 25284 19180 25396 19236
rect 25004 17726 25006 17778
rect 25058 17726 25060 17778
rect 22540 15428 22596 15438
rect 22428 15426 22596 15428
rect 22428 15374 22542 15426
rect 22594 15374 22596 15426
rect 22428 15372 22596 15374
rect 22540 15362 22596 15372
rect 21868 15262 21870 15314
rect 21922 15262 21924 15314
rect 21868 15250 21924 15262
rect 21420 14868 21476 14878
rect 21420 14642 21476 14812
rect 21420 14590 21422 14642
rect 21474 14590 21476 14642
rect 21420 14578 21476 14590
rect 22204 14530 22260 14542
rect 22204 14478 22206 14530
rect 22258 14478 22260 14530
rect 22204 13972 22260 14478
rect 22764 14532 22820 14542
rect 22764 14438 22820 14476
rect 22204 13906 22260 13916
rect 21308 13346 21364 13356
rect 21868 13412 21924 13422
rect 21084 13132 21812 13188
rect 21196 12964 21252 12974
rect 21532 12964 21588 12974
rect 21196 12870 21252 12908
rect 21308 12962 21588 12964
rect 21308 12910 21534 12962
rect 21586 12910 21588 12962
rect 21308 12908 21588 12910
rect 21308 12516 21364 12908
rect 21532 12898 21588 12908
rect 20524 12460 21364 12516
rect 21420 12738 21476 12750
rect 21420 12686 21422 12738
rect 21474 12686 21476 12738
rect 20524 12402 20580 12460
rect 20524 12350 20526 12402
rect 20578 12350 20580 12402
rect 20524 12338 20580 12350
rect 20300 12226 20356 12236
rect 20636 12292 20692 12302
rect 20636 12198 20692 12236
rect 20076 12178 20132 12190
rect 20076 12126 20078 12178
rect 20130 12126 20132 12178
rect 19852 11620 19908 11630
rect 19516 11618 19908 11620
rect 19516 11566 19854 11618
rect 19906 11566 19908 11618
rect 19516 11564 19908 11566
rect 19852 11554 19908 11564
rect 18956 11230 18958 11282
rect 19010 11230 19012 11282
rect 18956 11218 19012 11230
rect 20076 11284 20132 12126
rect 20412 12178 20468 12190
rect 20412 12126 20414 12178
rect 20466 12126 20468 12178
rect 20188 11508 20244 11518
rect 20188 11394 20244 11452
rect 20188 11342 20190 11394
rect 20242 11342 20244 11394
rect 20188 11330 20244 11342
rect 20412 11394 20468 12126
rect 21084 12066 21140 12078
rect 21084 12014 21086 12066
rect 21138 12014 21140 12066
rect 20412 11342 20414 11394
rect 20466 11342 20468 11394
rect 20076 11218 20132 11228
rect 19292 11172 19348 11182
rect 19964 11172 20020 11182
rect 19292 11170 20020 11172
rect 19292 11118 19294 11170
rect 19346 11118 19966 11170
rect 20018 11118 20020 11170
rect 19292 11116 20020 11118
rect 19292 10052 19348 11116
rect 19964 11106 20020 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19292 9986 19348 9996
rect 19628 10722 19684 10734
rect 19628 10670 19630 10722
rect 19682 10670 19684 10722
rect 18620 9938 18788 9940
rect 18620 9886 18622 9938
rect 18674 9886 18788 9938
rect 18620 9884 18788 9886
rect 18620 9874 18676 9884
rect 18172 9650 18228 9660
rect 19068 9716 19124 9726
rect 19068 9622 19124 9660
rect 19180 9604 19236 9614
rect 18732 9156 18788 9166
rect 18956 9156 19012 9166
rect 18732 9154 18956 9156
rect 18732 9102 18734 9154
rect 18786 9102 18956 9154
rect 18732 9100 18956 9102
rect 18732 9090 18788 9100
rect 18956 9062 19012 9100
rect 19068 8930 19124 8942
rect 19068 8878 19070 8930
rect 19122 8878 19124 8930
rect 17052 8318 17054 8370
rect 17106 8318 17108 8370
rect 17052 8306 17108 8318
rect 18844 8484 18900 8494
rect 16380 8206 16382 8258
rect 16434 8206 16436 8258
rect 16380 8194 16436 8206
rect 16044 8148 16100 8158
rect 15036 8034 15092 8046
rect 15036 7982 15038 8034
rect 15090 7982 15092 8034
rect 15036 7812 15092 7982
rect 15036 7746 15092 7756
rect 14924 7634 14980 7644
rect 16044 7700 16100 8092
rect 13916 7586 14196 7588
rect 13916 7534 13918 7586
rect 13970 7534 14196 7586
rect 13916 7532 14196 7534
rect 13916 7522 13972 7532
rect 16044 7362 16100 7644
rect 16492 7476 16548 7486
rect 16492 7382 16548 7420
rect 16044 7310 16046 7362
rect 16098 7310 16100 7362
rect 16044 7298 16100 7310
rect 13356 6514 13412 6524
rect 1708 6468 1764 6478
rect 1708 6374 1764 6412
rect 1708 6018 1764 6030
rect 1708 5966 1710 6018
rect 1762 5966 1764 6018
rect 1708 5460 1764 5966
rect 18844 5906 18900 8428
rect 19068 8372 19124 8878
rect 19068 8306 19124 8316
rect 19180 8370 19236 9548
rect 19180 8318 19182 8370
rect 19234 8318 19236 8370
rect 19180 8306 19236 8318
rect 19292 9042 19348 9054
rect 19292 8990 19294 9042
rect 19346 8990 19348 9042
rect 19292 8148 19348 8990
rect 19292 8082 19348 8092
rect 19404 9042 19460 9054
rect 19404 8990 19406 9042
rect 19458 8990 19460 9042
rect 19404 8036 19460 8990
rect 19628 9044 19684 10670
rect 19964 10724 20020 10734
rect 20020 10668 20132 10724
rect 19964 10658 20020 10668
rect 19740 10052 19796 10062
rect 19740 9714 19796 9996
rect 20076 9828 20132 10668
rect 20412 10164 20468 11342
rect 20412 10098 20468 10108
rect 20524 11508 20580 11518
rect 20524 9938 20580 11452
rect 21084 11508 21140 12014
rect 21084 11442 21140 11452
rect 21308 11284 21364 11294
rect 21308 11190 21364 11228
rect 21420 10388 21476 12686
rect 20860 10332 21476 10388
rect 21532 11394 21588 11406
rect 21532 11342 21534 11394
rect 21586 11342 21588 11394
rect 20524 9886 20526 9938
rect 20578 9886 20580 9938
rect 20524 9828 20580 9886
rect 20748 9940 20804 9950
rect 20748 9846 20804 9884
rect 20076 9772 20244 9828
rect 19740 9662 19742 9714
rect 19794 9662 19796 9714
rect 19740 9650 19796 9662
rect 20076 9604 20132 9642
rect 20076 9538 20132 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20188 9268 20244 9772
rect 20524 9762 20580 9772
rect 20860 9380 20916 10332
rect 21420 10164 21476 10174
rect 21420 10050 21476 10108
rect 21420 9998 21422 10050
rect 21474 9998 21476 10050
rect 21420 9986 21476 9998
rect 21532 9940 21588 11342
rect 21756 10164 21812 13132
rect 21868 12962 21924 13356
rect 21868 12910 21870 12962
rect 21922 12910 21924 12962
rect 21868 12898 21924 12910
rect 23212 12404 23268 17388
rect 25004 16212 25060 17726
rect 25228 17780 25284 19180
rect 26012 19124 26068 19134
rect 25676 19122 26068 19124
rect 25676 19070 26014 19122
rect 26066 19070 26068 19122
rect 25676 19068 26068 19070
rect 25564 18562 25620 18574
rect 25564 18510 25566 18562
rect 25618 18510 25620 18562
rect 25340 18452 25396 18462
rect 25340 18358 25396 18396
rect 25564 18340 25620 18510
rect 25564 18274 25620 18284
rect 25676 18338 25732 19068
rect 26012 19058 26068 19068
rect 25676 18286 25678 18338
rect 25730 18286 25732 18338
rect 25676 18274 25732 18286
rect 25228 17714 25284 17724
rect 25564 17780 25620 17790
rect 25004 16146 25060 16156
rect 25564 16210 25620 17724
rect 25564 16158 25566 16210
rect 25618 16158 25620 16210
rect 25564 16146 25620 16158
rect 25116 16100 25172 16110
rect 25116 16006 25172 16044
rect 25676 16100 25732 16110
rect 23436 15988 23492 15998
rect 23436 15894 23492 15932
rect 24332 15988 24388 15998
rect 24332 15894 24388 15932
rect 24668 15986 24724 15998
rect 24668 15934 24670 15986
rect 24722 15934 24724 15986
rect 23324 15874 23380 15886
rect 23324 15822 23326 15874
rect 23378 15822 23380 15874
rect 23324 14532 23380 15822
rect 23884 15204 23940 15214
rect 23884 14642 23940 15148
rect 23884 14590 23886 14642
rect 23938 14590 23940 14642
rect 23884 14578 23940 14590
rect 24668 15202 24724 15934
rect 24668 15150 24670 15202
rect 24722 15150 24724 15202
rect 23324 14466 23380 14476
rect 23436 14530 23492 14542
rect 23436 14478 23438 14530
rect 23490 14478 23492 14530
rect 23436 14084 23492 14478
rect 23772 14532 23828 14542
rect 23772 14438 23828 14476
rect 23996 14532 24052 14542
rect 23996 14438 24052 14476
rect 23436 14018 23492 14028
rect 24668 13972 24724 15150
rect 24780 15988 24836 15998
rect 24780 14418 24836 15932
rect 25676 15426 25732 16044
rect 25676 15374 25678 15426
rect 25730 15374 25732 15426
rect 25676 15362 25732 15374
rect 25340 15204 25396 15242
rect 25340 15138 25396 15148
rect 26124 15148 26180 19852
rect 26236 19460 26292 20076
rect 26348 20018 26404 20030
rect 26348 19966 26350 20018
rect 26402 19966 26404 20018
rect 26348 19796 26404 19966
rect 26684 20020 26740 20030
rect 26684 19926 26740 19964
rect 26348 19730 26404 19740
rect 26460 19908 26516 19918
rect 26236 19394 26292 19404
rect 26348 18564 26404 18574
rect 26460 18564 26516 19852
rect 26348 18562 26516 18564
rect 26348 18510 26350 18562
rect 26402 18510 26516 18562
rect 26348 18508 26516 18510
rect 26572 19460 26628 19470
rect 26348 18498 26404 18508
rect 26572 18450 26628 19404
rect 26572 18398 26574 18450
rect 26626 18398 26628 18450
rect 26572 18386 26628 18398
rect 26684 18452 26740 18462
rect 26684 17444 26740 18396
rect 26684 17350 26740 17388
rect 26124 15092 26516 15148
rect 25116 14532 25172 14542
rect 25900 14532 25956 14542
rect 25116 14438 25172 14476
rect 25676 14530 25956 14532
rect 25676 14478 25902 14530
rect 25954 14478 25956 14530
rect 25676 14476 25956 14478
rect 24780 14366 24782 14418
rect 24834 14366 24836 14418
rect 24780 14354 24836 14366
rect 24668 13906 24724 13916
rect 25340 14084 25396 14094
rect 25340 13970 25396 14028
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 25452 13972 25508 13982
rect 25452 13878 25508 13916
rect 25676 13858 25732 14476
rect 25900 14466 25956 14476
rect 25900 14308 25956 14318
rect 25676 13806 25678 13858
rect 25730 13806 25732 13858
rect 25228 13746 25284 13758
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 25228 13188 25284 13694
rect 25228 13122 25284 13132
rect 25564 12852 25620 12862
rect 25452 12850 25620 12852
rect 25452 12798 25566 12850
rect 25618 12798 25620 12850
rect 25452 12796 25620 12798
rect 25452 12404 25508 12796
rect 25564 12786 25620 12796
rect 23212 11508 23268 12348
rect 25116 12402 25508 12404
rect 25116 12350 25454 12402
rect 25506 12350 25508 12402
rect 25116 12348 25508 12350
rect 22988 11506 23268 11508
rect 22988 11454 23214 11506
rect 23266 11454 23268 11506
rect 22988 11452 23268 11454
rect 22988 10610 23044 11452
rect 23212 11442 23268 11452
rect 24332 11956 24388 11966
rect 24332 10722 24388 11900
rect 24444 11844 24500 11854
rect 24444 11394 24500 11788
rect 25116 11506 25172 12348
rect 25452 12338 25508 12348
rect 25228 11956 25284 11966
rect 25228 11862 25284 11900
rect 25564 11956 25620 11966
rect 25564 11862 25620 11900
rect 25116 11454 25118 11506
rect 25170 11454 25172 11506
rect 25116 11442 25172 11454
rect 24444 11342 24446 11394
rect 24498 11342 24500 11394
rect 24444 11330 24500 11342
rect 25004 11396 25060 11406
rect 24332 10670 24334 10722
rect 24386 10670 24388 10722
rect 24332 10658 24388 10670
rect 22988 10558 22990 10610
rect 23042 10558 23044 10610
rect 22988 10546 23044 10558
rect 23660 10610 23716 10622
rect 23660 10558 23662 10610
rect 23714 10558 23716 10610
rect 21532 9874 21588 9884
rect 21644 10108 21812 10164
rect 21868 10164 21924 10174
rect 21308 9716 21364 9726
rect 21308 9622 21364 9660
rect 20076 9212 20244 9268
rect 20636 9324 20916 9380
rect 19852 9044 19908 9054
rect 19628 9042 19908 9044
rect 19628 8990 19854 9042
rect 19906 8990 19908 9042
rect 19628 8988 19908 8990
rect 19852 8484 19908 8988
rect 19852 8418 19908 8428
rect 20076 8370 20132 9212
rect 20636 9154 20692 9324
rect 20636 9102 20638 9154
rect 20690 9102 20692 9154
rect 20636 9090 20692 9102
rect 21644 8484 21700 10108
rect 21868 10052 21924 10108
rect 23660 10164 23716 10558
rect 23660 10098 23716 10108
rect 24220 10610 24276 10622
rect 24220 10558 24222 10610
rect 24274 10558 24276 10610
rect 21756 9996 21924 10052
rect 21756 9826 21812 9996
rect 22316 9938 22372 9950
rect 22316 9886 22318 9938
rect 22370 9886 22372 9938
rect 21756 9774 21758 9826
rect 21810 9774 21812 9826
rect 21756 9762 21812 9774
rect 22204 9828 22260 9838
rect 22316 9828 22372 9886
rect 23436 9940 23492 9950
rect 23212 9828 23268 9838
rect 22316 9826 23268 9828
rect 22316 9774 23214 9826
rect 23266 9774 23268 9826
rect 22316 9772 23268 9774
rect 21084 8428 21700 8484
rect 20076 8318 20078 8370
rect 20130 8318 20132 8370
rect 19964 8260 20020 8270
rect 19404 7970 19460 7980
rect 19516 8258 20020 8260
rect 19516 8206 19966 8258
rect 20018 8206 20020 8258
rect 19516 8204 20020 8206
rect 19516 6018 19572 8204
rect 19964 8194 20020 8204
rect 19740 8036 19796 8046
rect 20076 8036 20132 8318
rect 20300 8372 20356 8382
rect 20300 8278 20356 8316
rect 20524 8260 20580 8270
rect 20524 8166 20580 8204
rect 19740 8034 20132 8036
rect 19740 7982 19742 8034
rect 19794 7982 20132 8034
rect 19740 7980 20132 7982
rect 19740 7970 19796 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 21084 7698 21140 8428
rect 21084 7646 21086 7698
rect 21138 7646 21140 7698
rect 21084 7634 21140 7646
rect 21308 8260 21364 8270
rect 21308 6690 21364 8204
rect 21644 8258 21700 8428
rect 21644 8206 21646 8258
rect 21698 8206 21700 8258
rect 21644 8194 21700 8206
rect 21980 9602 22036 9614
rect 21980 9550 21982 9602
rect 22034 9550 22036 9602
rect 21420 8146 21476 8158
rect 21420 8094 21422 8146
rect 21474 8094 21476 8146
rect 21420 8036 21476 8094
rect 21532 8148 21588 8158
rect 21532 8054 21588 8092
rect 21420 7970 21476 7980
rect 21644 7812 21700 7822
rect 21308 6638 21310 6690
rect 21362 6638 21364 6690
rect 21308 6626 21364 6638
rect 21532 6692 21588 6702
rect 21532 6598 21588 6636
rect 21420 6466 21476 6478
rect 21420 6414 21422 6466
rect 21474 6414 21476 6466
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19516 5966 19518 6018
rect 19570 5966 19572 6018
rect 19516 5954 19572 5966
rect 18844 5854 18846 5906
rect 18898 5854 18900 5906
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 1708 5394 1764 5404
rect 18844 5124 18900 5854
rect 21308 5348 21364 5358
rect 21420 5348 21476 6414
rect 21644 5794 21700 7756
rect 21980 7812 22036 9550
rect 22204 9380 22260 9772
rect 23212 9762 23268 9772
rect 23436 9826 23492 9884
rect 23660 9940 23716 9950
rect 23660 9846 23716 9884
rect 23436 9774 23438 9826
rect 23490 9774 23492 9826
rect 23436 9762 23492 9774
rect 23884 9826 23940 9838
rect 23884 9774 23886 9826
rect 23938 9774 23940 9826
rect 22204 9314 22260 9324
rect 22316 9602 22372 9614
rect 22316 9550 22318 9602
rect 22370 9550 22372 9602
rect 22092 8260 22148 8270
rect 22148 8204 22260 8260
rect 22092 8166 22148 8204
rect 21980 7746 22036 7756
rect 21868 6690 21924 6702
rect 21868 6638 21870 6690
rect 21922 6638 21924 6690
rect 21868 6580 21924 6638
rect 21868 6514 21924 6524
rect 21980 6692 22036 6702
rect 21980 5906 22036 6636
rect 21980 5854 21982 5906
rect 22034 5854 22036 5906
rect 21980 5842 22036 5854
rect 22204 5906 22260 8204
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 22204 5842 22260 5854
rect 22316 6690 22372 9550
rect 22764 9604 22820 9614
rect 22540 9268 22596 9278
rect 22428 8034 22484 8046
rect 22428 7982 22430 8034
rect 22482 7982 22484 8034
rect 22428 7812 22484 7982
rect 22428 7746 22484 7756
rect 22316 6638 22318 6690
rect 22370 6638 22372 6690
rect 21644 5742 21646 5794
rect 21698 5742 21700 5794
rect 21644 5730 21700 5742
rect 21308 5346 21476 5348
rect 21308 5294 21310 5346
rect 21362 5294 21476 5346
rect 21308 5292 21476 5294
rect 21644 5348 21700 5358
rect 21308 5282 21364 5292
rect 18844 5058 18900 5068
rect 19516 5124 19572 5134
rect 1708 4900 1764 4910
rect 1708 4806 1764 4844
rect 1708 4450 1764 4462
rect 1708 4398 1710 4450
rect 1762 4398 1764 4450
rect 1708 4116 1764 4398
rect 19516 4338 19572 5068
rect 21644 5122 21700 5292
rect 21644 5070 21646 5122
rect 21698 5070 21700 5122
rect 21644 5058 21700 5070
rect 21420 4898 21476 4910
rect 21420 4846 21422 4898
rect 21474 4846 21476 4898
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 21420 4676 21476 4846
rect 19836 4666 20100 4676
rect 20188 4620 21476 4676
rect 19516 4286 19518 4338
rect 19570 4286 19572 4338
rect 19516 4274 19572 4286
rect 19852 4564 19908 4574
rect 1708 4050 1764 4060
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 19516 3668 19572 3678
rect 1708 3444 1764 3454
rect 1708 3330 1764 3388
rect 10332 3332 10388 3342
rect 11004 3332 11060 3342
rect 1708 3278 1710 3330
rect 1762 3278 1764 3330
rect 1708 3266 1764 3278
rect 10108 3330 10388 3332
rect 10108 3278 10334 3330
rect 10386 3278 10388 3330
rect 10108 3276 10388 3278
rect 10108 800 10164 3276
rect 10332 3266 10388 3276
rect 10780 3330 11060 3332
rect 10780 3278 11006 3330
rect 11058 3278 11060 3330
rect 10780 3276 11060 3278
rect 10780 800 10836 3276
rect 11004 3266 11060 3276
rect 19516 800 19572 3612
rect 19628 3444 19684 3482
rect 19628 3378 19684 3388
rect 19852 3442 19908 4508
rect 20188 4450 20244 4620
rect 20188 4398 20190 4450
rect 20242 4398 20244 4450
rect 20188 4386 20244 4398
rect 22316 4226 22372 6638
rect 22540 6692 22596 9212
rect 22764 8930 22820 9548
rect 22876 9602 22932 9614
rect 22876 9550 22878 9602
rect 22930 9550 22932 9602
rect 22876 9380 22932 9550
rect 22876 9314 22932 9324
rect 23772 9268 23828 9278
rect 23772 9154 23828 9212
rect 23772 9102 23774 9154
rect 23826 9102 23828 9154
rect 23772 9090 23828 9102
rect 23884 9156 23940 9774
rect 23884 9062 23940 9100
rect 24220 9826 24276 10558
rect 24220 9774 24222 9826
rect 24274 9774 24276 9826
rect 22764 8878 22766 8930
rect 22818 8878 22820 8930
rect 22764 8866 22820 8878
rect 22764 8148 22820 8158
rect 22764 8054 22820 8092
rect 24220 8148 24276 9774
rect 24556 10612 24612 10622
rect 24444 9604 24500 9614
rect 24444 9510 24500 9548
rect 24332 9492 24388 9502
rect 24332 9042 24388 9436
rect 24556 9266 24612 10556
rect 25004 10276 25060 11340
rect 25452 10836 25508 10846
rect 25676 10836 25732 13806
rect 25452 10834 25732 10836
rect 25452 10782 25454 10834
rect 25506 10782 25732 10834
rect 25452 10780 25732 10782
rect 25788 14252 25900 14308
rect 25452 10770 25508 10780
rect 25340 10612 25396 10622
rect 25340 10518 25396 10556
rect 25564 10610 25620 10622
rect 25564 10558 25566 10610
rect 25618 10558 25620 10610
rect 25004 10220 25396 10276
rect 24780 9940 24836 9950
rect 24780 9938 25172 9940
rect 24780 9886 24782 9938
rect 24834 9886 25172 9938
rect 24780 9884 25172 9886
rect 24780 9874 24836 9884
rect 24780 9716 24836 9726
rect 24780 9622 24836 9660
rect 24556 9214 24558 9266
rect 24610 9214 24612 9266
rect 24556 9202 24612 9214
rect 24668 9602 24724 9614
rect 24668 9550 24670 9602
rect 24722 9550 24724 9602
rect 24668 9268 24724 9550
rect 24668 9202 24724 9212
rect 25116 9156 25172 9884
rect 25340 9938 25396 10220
rect 25340 9886 25342 9938
rect 25394 9886 25396 9938
rect 25340 9874 25396 9886
rect 25564 9940 25620 10558
rect 25564 9874 25620 9884
rect 25228 9604 25284 9614
rect 25228 9510 25284 9548
rect 25676 9268 25732 9278
rect 25676 9174 25732 9212
rect 25228 9156 25284 9166
rect 25116 9154 25284 9156
rect 25116 9102 25230 9154
rect 25282 9102 25284 9154
rect 25116 9100 25284 9102
rect 25228 9090 25284 9100
rect 25452 9156 25508 9166
rect 25452 9062 25508 9100
rect 24332 8990 24334 9042
rect 24386 8990 24388 9042
rect 24332 8978 24388 8990
rect 24668 9044 24724 9054
rect 24668 8950 24724 8988
rect 24220 8082 24276 8092
rect 25788 7924 25844 14252
rect 25900 14242 25956 14252
rect 26012 13524 26068 13534
rect 26012 12850 26068 13468
rect 26012 12798 26014 12850
rect 26066 12798 26068 12850
rect 26012 12786 26068 12798
rect 26348 12962 26404 12974
rect 26348 12910 26350 12962
rect 26402 12910 26404 12962
rect 26348 11956 26404 12910
rect 26348 11890 26404 11900
rect 26012 10610 26068 10622
rect 26012 10558 26014 10610
rect 26066 10558 26068 10610
rect 25900 9828 25956 9838
rect 25900 9044 25956 9772
rect 26012 9266 26068 10558
rect 26012 9214 26014 9266
rect 26066 9214 26068 9266
rect 26012 9202 26068 9214
rect 26236 10052 26292 10062
rect 26236 9380 26292 9996
rect 26348 9940 26404 9950
rect 26348 9714 26404 9884
rect 26348 9662 26350 9714
rect 26402 9662 26404 9714
rect 26348 9650 26404 9662
rect 26236 9266 26292 9324
rect 26236 9214 26238 9266
rect 26290 9214 26292 9266
rect 26236 9202 26292 9214
rect 26348 9044 26404 9054
rect 25900 9042 26180 9044
rect 25900 8990 25902 9042
rect 25954 8990 26180 9042
rect 25900 8988 26180 8990
rect 25900 8978 25956 8988
rect 26124 8370 26180 8988
rect 26124 8318 26126 8370
rect 26178 8318 26180 8370
rect 26124 8306 26180 8318
rect 25340 7868 25844 7924
rect 26348 8036 26404 8988
rect 25228 6804 25284 6814
rect 22540 6578 22596 6636
rect 24668 6802 25284 6804
rect 24668 6750 25230 6802
rect 25282 6750 25284 6802
rect 24668 6748 25284 6750
rect 22540 6526 22542 6578
rect 22594 6526 22596 6578
rect 22540 6514 22596 6526
rect 22988 6580 23044 6590
rect 22988 6486 23044 6524
rect 24220 6578 24276 6590
rect 24220 6526 24222 6578
rect 24274 6526 24276 6578
rect 24108 6468 24164 6478
rect 23212 6132 23268 6142
rect 23212 6038 23268 6076
rect 23436 6020 23492 6030
rect 23436 5926 23492 5964
rect 23100 5906 23156 5918
rect 23100 5854 23102 5906
rect 23154 5854 23156 5906
rect 22540 5684 22596 5694
rect 23100 5684 23156 5854
rect 24108 5906 24164 6412
rect 24108 5854 24110 5906
rect 24162 5854 24164 5906
rect 24108 5842 24164 5854
rect 24220 6020 24276 6526
rect 24332 6580 24388 6590
rect 24332 6486 24388 6524
rect 24556 6468 24612 6478
rect 24220 5794 24276 5964
rect 24220 5742 24222 5794
rect 24274 5742 24276 5794
rect 24220 5730 24276 5742
rect 24444 6466 24612 6468
rect 24444 6414 24558 6466
rect 24610 6414 24612 6466
rect 24444 6412 24612 6414
rect 22540 5682 23156 5684
rect 22540 5630 22542 5682
rect 22594 5630 23156 5682
rect 22540 5628 23156 5630
rect 22540 5618 22596 5628
rect 23100 5348 23156 5628
rect 23100 5282 23156 5292
rect 22876 5124 22932 5134
rect 22876 5030 22932 5068
rect 24108 5124 24164 5134
rect 23660 5012 23716 5022
rect 23660 5010 24052 5012
rect 23660 4958 23662 5010
rect 23714 4958 24052 5010
rect 23660 4956 24052 4958
rect 23660 4946 23716 4956
rect 22316 4174 22318 4226
rect 22370 4174 22372 4226
rect 22316 4162 22372 4174
rect 23996 4226 24052 4956
rect 24108 4562 24164 5068
rect 24108 4510 24110 4562
rect 24162 4510 24164 4562
rect 24108 4498 24164 4510
rect 24332 4452 24388 4462
rect 24444 4452 24500 6412
rect 24556 6402 24612 6412
rect 24668 6018 24724 6748
rect 25228 6738 25284 6748
rect 24892 6580 24948 6590
rect 25340 6580 25396 7868
rect 24948 6524 25396 6580
rect 25452 7700 25508 7710
rect 25452 6804 25508 7644
rect 25564 6916 25620 6926
rect 25564 6914 26292 6916
rect 25564 6862 25566 6914
rect 25618 6862 26292 6914
rect 25564 6860 26292 6862
rect 25564 6850 25620 6860
rect 25452 6578 25508 6748
rect 25452 6526 25454 6578
rect 25506 6526 25508 6578
rect 24892 6486 24948 6524
rect 25452 6514 25508 6526
rect 26012 6578 26068 6590
rect 26012 6526 26014 6578
rect 26066 6526 26068 6578
rect 25900 6466 25956 6478
rect 25900 6414 25902 6466
rect 25954 6414 25956 6466
rect 25900 6356 25956 6414
rect 25900 6290 25956 6300
rect 26012 6132 26068 6526
rect 24668 5966 24670 6018
rect 24722 5966 24724 6018
rect 24668 5954 24724 5966
rect 25788 6076 26012 6132
rect 25564 5908 25620 5918
rect 25564 5814 25620 5852
rect 25788 5236 25844 6076
rect 26012 6066 26068 6076
rect 26236 6018 26292 6860
rect 26348 6356 26404 7980
rect 26460 6804 26516 15092
rect 26572 14418 26628 14430
rect 26572 14366 26574 14418
rect 26626 14366 26628 14418
rect 26572 14084 26628 14366
rect 26796 14308 26852 21420
rect 27580 20132 27636 20142
rect 27692 20132 27748 21422
rect 28140 20804 28196 21646
rect 28140 20738 28196 20748
rect 27580 20130 27748 20132
rect 27580 20078 27582 20130
rect 27634 20078 27748 20130
rect 27580 20076 27748 20078
rect 27580 20066 27636 20076
rect 27020 20020 27076 20030
rect 27020 19684 27076 19964
rect 27244 20020 27300 20030
rect 27244 19926 27300 19964
rect 27468 19908 27524 19918
rect 27468 19814 27524 19852
rect 27020 19618 27076 19628
rect 27244 18452 27300 18462
rect 27244 18358 27300 18396
rect 26908 18226 26964 18238
rect 26908 18174 26910 18226
rect 26962 18174 26964 18226
rect 26908 17780 26964 18174
rect 27020 17780 27076 17790
rect 27468 17780 27524 17790
rect 26908 17778 27524 17780
rect 26908 17726 27022 17778
rect 27074 17726 27470 17778
rect 27522 17726 27524 17778
rect 26908 17724 27524 17726
rect 27020 17714 27076 17724
rect 27468 17714 27524 17724
rect 27692 17666 27748 20076
rect 28364 20020 28420 22428
rect 28476 22260 28532 22270
rect 28476 22166 28532 22204
rect 28588 21028 28644 26012
rect 28700 21140 28756 26852
rect 29484 26852 29540 26862
rect 29484 26758 29540 26796
rect 29596 26852 29764 26908
rect 29932 26964 29988 26974
rect 29484 25396 29540 25406
rect 29372 25394 29540 25396
rect 29372 25342 29486 25394
rect 29538 25342 29540 25394
rect 29372 25340 29540 25342
rect 29148 23268 29204 23278
rect 28924 23212 29148 23268
rect 28924 21810 28980 23212
rect 29148 23202 29204 23212
rect 29036 22596 29092 22606
rect 29036 22502 29092 22540
rect 29372 22372 29428 25340
rect 29484 25330 29540 25340
rect 29484 23044 29540 23054
rect 29596 23044 29652 26852
rect 29708 25396 29764 25406
rect 29932 25396 29988 26908
rect 30492 26178 30548 26190
rect 30492 26126 30494 26178
rect 30546 26126 30548 26178
rect 30268 25508 30324 25518
rect 30492 25508 30548 26126
rect 30716 26066 30772 29932
rect 30828 29922 30884 29932
rect 31164 29986 31220 30492
rect 31276 30322 31332 32508
rect 31388 32562 31444 32732
rect 31388 32510 31390 32562
rect 31442 32510 31444 32562
rect 31388 32228 31444 32510
rect 31388 32162 31444 32172
rect 31500 32564 31556 33068
rect 31612 33122 31668 33180
rect 31612 33070 31614 33122
rect 31666 33070 31668 33122
rect 31612 32676 31668 33070
rect 31612 32610 31668 32620
rect 31500 32450 31556 32508
rect 31500 32398 31502 32450
rect 31554 32398 31556 32450
rect 31388 31780 31444 31790
rect 31500 31780 31556 32398
rect 31388 31778 31556 31780
rect 31388 31726 31390 31778
rect 31442 31726 31556 31778
rect 31388 31724 31556 31726
rect 31724 31780 31780 37212
rect 31836 35812 31892 37774
rect 32172 37828 32228 37838
rect 32172 37734 32228 37772
rect 31836 35746 31892 35756
rect 32060 37380 32116 37390
rect 31836 34018 31892 34030
rect 31836 33966 31838 34018
rect 31890 33966 31892 34018
rect 31836 33906 31892 33966
rect 31836 33854 31838 33906
rect 31890 33854 31892 33906
rect 31836 33842 31892 33854
rect 32060 33124 32116 37324
rect 32396 37044 32452 38780
rect 32508 37828 32564 37838
rect 32508 37268 32564 37772
rect 32508 37202 32564 37212
rect 32396 36978 32452 36988
rect 32284 35812 32340 35822
rect 32284 35718 32340 35756
rect 32508 35700 32564 35710
rect 32508 35606 32564 35644
rect 32172 35586 32228 35598
rect 32172 35534 32174 35586
rect 32226 35534 32228 35586
rect 32172 35476 32228 35534
rect 32172 35410 32228 35420
rect 32396 34802 32452 34814
rect 32396 34750 32398 34802
rect 32450 34750 32452 34802
rect 32396 34356 32452 34750
rect 32396 34290 32452 34300
rect 32284 34132 32340 34142
rect 32284 34038 32340 34076
rect 32172 33572 32228 33582
rect 32172 33478 32228 33516
rect 32284 33460 32340 33470
rect 32284 33234 32340 33404
rect 32284 33182 32286 33234
rect 32338 33182 32340 33234
rect 32172 33124 32228 33134
rect 32060 33122 32228 33124
rect 32060 33070 32174 33122
rect 32226 33070 32228 33122
rect 32060 33068 32228 33070
rect 31836 32900 31892 32910
rect 31836 32674 31892 32844
rect 32172 32788 32228 33068
rect 32172 32722 32228 32732
rect 31836 32622 31838 32674
rect 31890 32622 31892 32674
rect 31836 32610 31892 32622
rect 31836 31780 31892 31790
rect 31724 31724 31836 31780
rect 31388 31714 31444 31724
rect 31276 30270 31278 30322
rect 31330 30270 31332 30322
rect 31276 30258 31332 30270
rect 31836 30210 31892 31724
rect 32060 30324 32116 30334
rect 32284 30324 32340 33182
rect 32396 30324 32452 30334
rect 32284 30322 32452 30324
rect 32284 30270 32398 30322
rect 32450 30270 32452 30322
rect 32284 30268 32452 30270
rect 32060 30230 32116 30268
rect 31836 30158 31838 30210
rect 31890 30158 31892 30210
rect 31836 30146 31892 30158
rect 32172 30212 32228 30222
rect 32172 30098 32228 30156
rect 32172 30046 32174 30098
rect 32226 30046 32228 30098
rect 31164 29934 31166 29986
rect 31218 29934 31220 29986
rect 30828 29428 30884 29438
rect 30828 29334 30884 29372
rect 30940 28756 30996 28766
rect 30940 26292 30996 28700
rect 31164 27412 31220 29934
rect 31388 29986 31444 29998
rect 31388 29934 31390 29986
rect 31442 29934 31444 29986
rect 31388 29428 31444 29934
rect 31836 29876 31892 29886
rect 31836 29538 31892 29820
rect 31948 29764 32004 29774
rect 31948 29650 32004 29708
rect 31948 29598 31950 29650
rect 32002 29598 32004 29650
rect 31948 29586 32004 29598
rect 31836 29486 31838 29538
rect 31890 29486 31892 29538
rect 31836 29474 31892 29486
rect 31500 29428 31556 29438
rect 31388 29372 31500 29428
rect 31500 28754 31556 29372
rect 31500 28702 31502 28754
rect 31554 28702 31556 28754
rect 31500 28690 31556 28702
rect 31276 28644 31332 28654
rect 31276 28550 31332 28588
rect 32172 28644 32228 30046
rect 32396 29652 32452 30268
rect 32732 30212 32788 38892
rect 33068 38946 33124 39564
rect 40124 39396 40180 39406
rect 40124 39394 40292 39396
rect 40124 39342 40126 39394
rect 40178 39342 40292 39394
rect 40124 39340 40292 39342
rect 40124 39330 40180 39340
rect 40236 39060 40292 39340
rect 40348 39060 40404 39070
rect 40236 39004 40348 39060
rect 40348 38994 40404 39004
rect 33068 38894 33070 38946
rect 33122 38894 33124 38946
rect 33068 38882 33124 38894
rect 33292 38946 33348 38958
rect 33292 38894 33294 38946
rect 33346 38894 33348 38946
rect 33180 38724 33236 38734
rect 33180 38630 33236 38668
rect 33292 37828 33348 38894
rect 40124 38946 40180 38958
rect 40124 38894 40126 38946
rect 40178 38894 40180 38946
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 40124 38388 40180 38894
rect 40124 38322 40180 38332
rect 33292 37762 33348 37772
rect 40124 37826 40180 37838
rect 40124 37774 40126 37826
rect 40178 37774 40180 37826
rect 40124 37716 40180 37774
rect 40124 37650 40180 37660
rect 40124 37378 40180 37390
rect 40124 37326 40126 37378
rect 40178 37326 40180 37378
rect 32732 30146 32788 30156
rect 32844 37044 32900 37054
rect 32396 29586 32452 29596
rect 32620 29986 32676 29998
rect 32620 29934 32622 29986
rect 32674 29934 32676 29986
rect 32620 29428 32676 29934
rect 32844 29986 32900 36988
rect 40124 37044 40180 37326
rect 40124 36978 40180 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 33068 35700 33124 35710
rect 33068 35606 33124 35644
rect 33180 35586 33236 35598
rect 33180 35534 33182 35586
rect 33234 35534 33236 35586
rect 33068 34244 33124 34254
rect 33180 34244 33236 35534
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34524 35028 34580 35038
rect 33068 34242 33236 34244
rect 33068 34190 33070 34242
rect 33122 34190 33236 34242
rect 33068 34188 33236 34190
rect 33964 35026 34580 35028
rect 33964 34974 34526 35026
rect 34578 34974 34580 35026
rect 33964 34972 34580 34974
rect 33068 34178 33124 34188
rect 33516 34130 33572 34142
rect 33516 34078 33518 34130
rect 33570 34078 33572 34130
rect 33516 33348 33572 34078
rect 33964 34132 34020 34972
rect 34524 34962 34580 34972
rect 33964 34130 34132 34132
rect 33964 34078 33966 34130
rect 34018 34078 34132 34130
rect 33964 34076 34132 34078
rect 33964 34066 34020 34076
rect 33292 33292 33516 33348
rect 33292 32786 33348 33292
rect 33516 33282 33572 33292
rect 33292 32734 33294 32786
rect 33346 32734 33348 32786
rect 33292 32722 33348 32734
rect 33628 32674 33684 32686
rect 33628 32622 33630 32674
rect 33682 32622 33684 32674
rect 33404 32452 33460 32462
rect 33404 32228 33460 32396
rect 33628 32340 33684 32622
rect 33964 32452 34020 32462
rect 33964 32358 34020 32396
rect 33628 32274 33684 32284
rect 33292 32172 33460 32228
rect 33292 31666 33348 32172
rect 33404 31780 33460 31790
rect 33740 31780 33796 31790
rect 33404 31778 33796 31780
rect 33404 31726 33406 31778
rect 33458 31726 33742 31778
rect 33794 31726 33796 31778
rect 33404 31724 33796 31726
rect 33404 31714 33460 31724
rect 33740 31714 33796 31724
rect 33292 31614 33294 31666
rect 33346 31614 33348 31666
rect 33292 31602 33348 31614
rect 32956 30212 33012 30222
rect 32956 30118 33012 30156
rect 33964 30212 34020 30222
rect 34076 30212 34132 34076
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34412 33348 34468 33358
rect 34412 32562 34468 33292
rect 35196 33346 35252 33358
rect 35196 33294 35198 33346
rect 35250 33294 35252 33346
rect 34972 33236 35028 33246
rect 35196 33236 35252 33294
rect 36204 33292 36484 33348
rect 35028 33180 35252 33236
rect 35868 33236 35924 33246
rect 36204 33236 36260 33292
rect 35924 33234 36260 33236
rect 35924 33182 36206 33234
rect 36258 33182 36260 33234
rect 35924 33180 36260 33182
rect 34972 33142 35028 33180
rect 35868 33142 35924 33180
rect 36204 33170 36260 33180
rect 35644 33122 35700 33134
rect 35644 33070 35646 33122
rect 35698 33070 35700 33122
rect 35644 32900 35700 33070
rect 35756 33124 35812 33134
rect 35756 33030 35812 33068
rect 36316 33122 36372 33134
rect 36316 33070 36318 33122
rect 36370 33070 36372 33122
rect 36316 32900 36372 33070
rect 35644 32844 36372 32900
rect 34412 32510 34414 32562
rect 34466 32510 34468 32562
rect 34412 32498 34468 32510
rect 35980 32562 36036 32574
rect 35980 32510 35982 32562
rect 36034 32510 36036 32562
rect 34748 32450 34804 32462
rect 34748 32398 34750 32450
rect 34802 32398 34804 32450
rect 34020 30156 34132 30212
rect 34188 32340 34244 32350
rect 34188 31778 34244 32284
rect 34636 31892 34692 31902
rect 34188 31726 34190 31778
rect 34242 31726 34244 31778
rect 34188 31332 34244 31726
rect 33964 30118 34020 30156
rect 32844 29934 32846 29986
rect 32898 29934 32900 29986
rect 32844 29876 32900 29934
rect 32844 29810 32900 29820
rect 33628 29986 33684 29998
rect 33628 29934 33630 29986
rect 33682 29934 33684 29986
rect 33292 29764 33348 29774
rect 33068 29428 33124 29438
rect 32620 29426 33124 29428
rect 32620 29374 33070 29426
rect 33122 29374 33124 29426
rect 32620 29372 33124 29374
rect 32172 28578 32228 28588
rect 31164 27346 31220 27356
rect 31724 28530 31780 28542
rect 31724 28478 31726 28530
rect 31778 28478 31780 28530
rect 31612 27188 31668 27198
rect 31612 27094 31668 27132
rect 31500 27074 31556 27086
rect 31500 27022 31502 27074
rect 31554 27022 31556 27074
rect 31388 26964 31444 27002
rect 31388 26898 31444 26908
rect 31388 26516 31444 26526
rect 31500 26516 31556 27022
rect 31724 27076 31780 28478
rect 32284 27972 32340 27982
rect 32284 27878 32340 27916
rect 31724 27010 31780 27020
rect 31836 27858 31892 27870
rect 31836 27806 31838 27858
rect 31890 27806 31892 27858
rect 31388 26514 31556 26516
rect 31388 26462 31390 26514
rect 31442 26462 31556 26514
rect 31388 26460 31556 26462
rect 31388 26450 31444 26460
rect 31724 26292 31780 26302
rect 30940 26198 30996 26236
rect 31388 26290 31780 26292
rect 31388 26238 31726 26290
rect 31778 26238 31780 26290
rect 31388 26236 31780 26238
rect 30716 26014 30718 26066
rect 30770 26014 30772 26066
rect 30716 26002 30772 26014
rect 31276 26068 31332 26078
rect 31388 26068 31444 26236
rect 31724 26226 31780 26236
rect 31276 26066 31444 26068
rect 31276 26014 31278 26066
rect 31330 26014 31444 26066
rect 31276 26012 31444 26014
rect 31500 26068 31556 26078
rect 31276 26002 31332 26012
rect 31500 25974 31556 26012
rect 31164 25620 31220 25630
rect 31164 25526 31220 25564
rect 30324 25452 30548 25508
rect 30828 25508 30884 25518
rect 30268 25414 30324 25452
rect 29708 25394 29988 25396
rect 29708 25342 29710 25394
rect 29762 25342 29934 25394
rect 29986 25342 29988 25394
rect 29708 25340 29988 25342
rect 29708 25330 29764 25340
rect 29932 25330 29988 25340
rect 30828 24834 30884 25452
rect 30828 24782 30830 24834
rect 30882 24782 30884 24834
rect 30828 24770 30884 24782
rect 31052 25506 31108 25518
rect 31052 25454 31054 25506
rect 31106 25454 31108 25506
rect 29820 23716 29876 23726
rect 29484 23042 29652 23044
rect 29484 22990 29486 23042
rect 29538 22990 29652 23042
rect 29484 22988 29652 22990
rect 29708 23714 29876 23716
rect 29708 23662 29822 23714
rect 29874 23662 29876 23714
rect 29708 23660 29876 23662
rect 29484 22978 29540 22988
rect 29708 22820 29764 23660
rect 29820 23650 29876 23660
rect 30492 23380 30548 23390
rect 30044 23268 30100 23278
rect 30044 23174 30100 23212
rect 28924 21758 28926 21810
rect 28978 21758 28980 21810
rect 28924 21746 28980 21758
rect 29036 22370 29428 22372
rect 29036 22318 29374 22370
rect 29426 22318 29428 22370
rect 29036 22316 29428 22318
rect 28812 21588 28868 21598
rect 29036 21588 29092 22316
rect 29372 22306 29428 22316
rect 29484 22764 29764 22820
rect 29820 23154 29876 23166
rect 29820 23102 29822 23154
rect 29874 23102 29876 23154
rect 29148 22148 29204 22158
rect 29484 22148 29540 22764
rect 29820 22372 29876 23102
rect 30492 23154 30548 23324
rect 30492 23102 30494 23154
rect 30546 23102 30548 23154
rect 30492 23090 30548 23102
rect 29932 23044 29988 23054
rect 29932 22950 29988 22988
rect 29820 22316 29988 22372
rect 29596 22260 29652 22270
rect 29596 22258 29876 22260
rect 29596 22206 29598 22258
rect 29650 22206 29876 22258
rect 29596 22204 29876 22206
rect 29596 22194 29652 22204
rect 29148 22054 29204 22092
rect 29372 22092 29540 22148
rect 28868 21532 29092 21588
rect 28812 21494 28868 21532
rect 28700 21084 28980 21140
rect 28588 20972 28868 21028
rect 28364 19954 28420 19964
rect 28140 19796 28196 19806
rect 28140 19346 28196 19740
rect 28140 19294 28142 19346
rect 28194 19294 28196 19346
rect 28140 19282 28196 19294
rect 28700 19572 28756 19582
rect 28588 19236 28644 19246
rect 28588 19142 28644 19180
rect 27692 17614 27694 17666
rect 27746 17614 27748 17666
rect 27692 17602 27748 17614
rect 28252 17666 28308 17678
rect 28252 17614 28254 17666
rect 28306 17614 28308 17666
rect 27132 17556 27188 17566
rect 27132 17462 27188 17500
rect 27916 17554 27972 17566
rect 27916 17502 27918 17554
rect 27970 17502 27972 17554
rect 27916 16324 27972 17502
rect 27916 16258 27972 16268
rect 27244 15426 27300 15438
rect 27244 15374 27246 15426
rect 27298 15374 27300 15426
rect 27244 14644 27300 15374
rect 27244 14578 27300 14588
rect 27468 15202 27524 15214
rect 27468 15150 27470 15202
rect 27522 15150 27524 15202
rect 26796 14242 26852 14252
rect 27132 14532 27188 14542
rect 26572 14028 26908 14084
rect 26852 13870 26908 14028
rect 26852 13858 26964 13870
rect 26852 13806 26910 13858
rect 26962 13806 26964 13858
rect 26852 13804 26964 13806
rect 26908 13794 26964 13804
rect 26684 13636 26740 13646
rect 26684 13186 26740 13580
rect 26684 13134 26686 13186
rect 26738 13134 26740 13186
rect 26684 13122 26740 13134
rect 27132 12852 27188 14476
rect 27468 13746 27524 15150
rect 28140 13748 28196 13758
rect 27468 13694 27470 13746
rect 27522 13694 27524 13746
rect 27468 13524 27524 13694
rect 27468 13458 27524 13468
rect 27580 13746 28196 13748
rect 27580 13694 28142 13746
rect 28194 13694 28196 13746
rect 27580 13692 28196 13694
rect 27244 13188 27300 13198
rect 27244 13094 27300 13132
rect 27132 12850 27300 12852
rect 27132 12798 27134 12850
rect 27186 12798 27300 12850
rect 27132 12796 27300 12798
rect 27132 12786 27188 12796
rect 26908 9826 26964 9838
rect 26908 9774 26910 9826
rect 26962 9774 26964 9826
rect 26908 9268 26964 9774
rect 26908 9202 26964 9212
rect 27132 9380 27188 9390
rect 27132 9042 27188 9324
rect 27132 8990 27134 9042
rect 27186 8990 27188 9042
rect 27132 8978 27188 8990
rect 27244 8428 27300 12796
rect 27580 10834 27636 13692
rect 28140 13682 28196 13692
rect 28252 13636 28308 17614
rect 28476 17442 28532 17454
rect 28476 17390 28478 17442
rect 28530 17390 28532 17442
rect 28476 16996 28532 17390
rect 28476 16930 28532 16940
rect 28588 16324 28644 16334
rect 28588 13970 28644 16268
rect 28700 14868 28756 19516
rect 28700 14802 28756 14812
rect 28588 13918 28590 13970
rect 28642 13918 28644 13970
rect 28588 13906 28644 13918
rect 28812 13972 28868 20972
rect 28812 13906 28868 13916
rect 28252 13570 28308 13580
rect 28924 13300 28980 21084
rect 29148 20690 29204 20702
rect 29148 20638 29150 20690
rect 29202 20638 29204 20690
rect 29148 18004 29204 20638
rect 29260 20578 29316 20590
rect 29260 20526 29262 20578
rect 29314 20526 29316 20578
rect 29260 19460 29316 20526
rect 29260 19394 29316 19404
rect 29372 20132 29428 22092
rect 29596 21700 29652 21710
rect 29596 21606 29652 21644
rect 29484 21586 29540 21598
rect 29484 21534 29486 21586
rect 29538 21534 29540 21586
rect 29484 21028 29540 21534
rect 29596 21364 29652 21374
rect 29596 21270 29652 21308
rect 29820 21028 29876 22204
rect 29932 22148 29988 22316
rect 29932 22082 29988 22092
rect 29484 20972 29652 21028
rect 29484 20804 29540 20814
rect 29484 20710 29540 20748
rect 29260 19236 29316 19246
rect 29372 19236 29428 20076
rect 29596 20580 29652 20972
rect 29708 20804 29764 20814
rect 29820 20804 29876 20972
rect 29708 20802 29876 20804
rect 29708 20750 29710 20802
rect 29762 20750 29876 20802
rect 29708 20748 29876 20750
rect 30156 21474 30212 21486
rect 30156 21422 30158 21474
rect 30210 21422 30212 21474
rect 29708 20738 29764 20748
rect 30156 20580 30212 21422
rect 30828 21028 30884 21038
rect 30828 20934 30884 20972
rect 29596 20524 30212 20580
rect 29484 19572 29540 19582
rect 29596 19572 29652 20524
rect 29932 20020 29988 20030
rect 29932 19926 29988 19964
rect 30380 20020 30436 20030
rect 29540 19516 29652 19572
rect 29484 19506 29540 19516
rect 29316 19180 29428 19236
rect 30380 19234 30436 19964
rect 30380 19182 30382 19234
rect 30434 19182 30436 19234
rect 29260 18562 29316 19180
rect 30380 19170 30436 19182
rect 29260 18510 29262 18562
rect 29314 18510 29316 18562
rect 29260 18498 29316 18510
rect 29484 19122 29540 19134
rect 29484 19070 29486 19122
rect 29538 19070 29540 19122
rect 29148 17948 29316 18004
rect 29148 17668 29204 17678
rect 29148 17574 29204 17612
rect 29148 16996 29204 17006
rect 29148 16902 29204 16940
rect 29260 15540 29316 17948
rect 29484 17668 29540 19070
rect 30604 19124 30660 19134
rect 30604 19030 30660 19068
rect 29820 19010 29876 19022
rect 29820 18958 29822 19010
rect 29874 18958 29876 19010
rect 29820 18676 29876 18958
rect 29820 18610 29876 18620
rect 30940 19010 30996 19022
rect 30940 18958 30942 19010
rect 30994 18958 30996 19010
rect 30716 17668 30772 17678
rect 30940 17668 30996 18958
rect 29484 17602 29540 17612
rect 30604 17666 30996 17668
rect 30604 17614 30718 17666
rect 30770 17614 30996 17666
rect 30604 17612 30996 17614
rect 30156 17556 30212 17566
rect 30492 17556 30548 17566
rect 30156 17554 30492 17556
rect 30156 17502 30158 17554
rect 30210 17502 30492 17554
rect 30156 17500 30492 17502
rect 30156 17490 30212 17500
rect 30492 17462 30548 17500
rect 29484 17444 29540 17454
rect 29820 17444 29876 17454
rect 29484 17442 29764 17444
rect 29484 17390 29486 17442
rect 29538 17390 29764 17442
rect 29484 17388 29764 17390
rect 29484 17378 29540 17388
rect 29484 16994 29540 17006
rect 29484 16942 29486 16994
rect 29538 16942 29540 16994
rect 29484 15876 29540 16942
rect 29708 15988 29764 17388
rect 29820 17442 29988 17444
rect 29820 17390 29822 17442
rect 29874 17390 29988 17442
rect 29820 17388 29988 17390
rect 29820 17378 29876 17388
rect 29932 16996 29988 17388
rect 30604 17332 30660 17612
rect 30716 17602 30772 17612
rect 30380 17276 30660 17332
rect 30716 17444 30772 17454
rect 29932 16882 29988 16940
rect 29932 16830 29934 16882
rect 29986 16830 29988 16882
rect 29932 16818 29988 16830
rect 30156 16994 30212 17006
rect 30156 16942 30158 16994
rect 30210 16942 30212 16994
rect 30156 16212 30212 16942
rect 30156 16146 30212 16156
rect 29708 15932 30100 15988
rect 29484 15810 29540 15820
rect 29820 15540 29876 15550
rect 29260 15538 29876 15540
rect 29260 15486 29822 15538
rect 29874 15486 29876 15538
rect 29260 15484 29876 15486
rect 29820 15474 29876 15484
rect 29932 15426 29988 15438
rect 29932 15374 29934 15426
rect 29986 15374 29988 15426
rect 29932 15092 29988 15374
rect 30044 15204 30100 15932
rect 30044 15138 30100 15148
rect 30156 15314 30212 15326
rect 30156 15262 30158 15314
rect 30210 15262 30212 15314
rect 29932 15026 29988 15036
rect 30156 15092 30212 15262
rect 30156 15026 30212 15036
rect 29820 14756 29876 14766
rect 29148 14644 29204 14654
rect 29148 14550 29204 14588
rect 29820 14530 29876 14700
rect 29820 14478 29822 14530
rect 29874 14478 29876 14530
rect 29820 14466 29876 14478
rect 30044 14530 30100 14542
rect 30044 14478 30046 14530
rect 30098 14478 30100 14530
rect 29820 13972 29876 13982
rect 29820 13878 29876 13916
rect 28924 13234 28980 13244
rect 27916 13188 27972 13198
rect 27916 12402 27972 13132
rect 29932 12740 29988 12750
rect 27916 12350 27918 12402
rect 27970 12350 27972 12402
rect 27916 12338 27972 12350
rect 29820 12738 29988 12740
rect 29820 12686 29934 12738
rect 29986 12686 29988 12738
rect 29820 12684 29988 12686
rect 28028 12180 28084 12190
rect 28028 12086 28084 12124
rect 28588 12180 28644 12190
rect 28588 12086 28644 12124
rect 29820 12180 29876 12684
rect 29932 12674 29988 12684
rect 30044 12516 30100 14478
rect 30156 13972 30212 13982
rect 30156 13858 30212 13916
rect 30156 13806 30158 13858
rect 30210 13806 30212 13858
rect 30156 12628 30212 13806
rect 30380 13860 30436 17276
rect 30492 16996 30548 17006
rect 30492 16902 30548 16940
rect 30492 15314 30548 15326
rect 30492 15262 30494 15314
rect 30546 15262 30548 15314
rect 30492 15148 30548 15262
rect 30716 15148 30772 17388
rect 30828 16994 30884 17006
rect 30828 16942 30830 16994
rect 30882 16942 30884 16994
rect 30828 16100 30884 16942
rect 30828 16034 30884 16044
rect 30940 15314 30996 15326
rect 30940 15262 30942 15314
rect 30994 15262 30996 15314
rect 30492 15092 30660 15148
rect 30716 15092 30884 15148
rect 30380 13794 30436 13804
rect 30492 14868 30548 14878
rect 30492 13970 30548 14812
rect 30492 13918 30494 13970
rect 30546 13918 30548 13970
rect 30492 13748 30548 13918
rect 30604 13972 30660 15092
rect 30828 14644 30884 15092
rect 30940 14868 30996 15262
rect 31052 15316 31108 25454
rect 31612 25396 31668 25406
rect 31612 25302 31668 25340
rect 31836 24946 31892 27806
rect 32060 27860 32116 27870
rect 32956 27860 33012 29372
rect 33068 29362 33124 29372
rect 33292 29426 33348 29708
rect 33292 29374 33294 29426
rect 33346 29374 33348 29426
rect 33292 29362 33348 29374
rect 33628 29428 33684 29934
rect 33628 29362 33684 29372
rect 34076 29876 34132 29886
rect 33852 29314 33908 29326
rect 33852 29262 33854 29314
rect 33906 29262 33908 29314
rect 33852 29204 33908 29262
rect 33404 29148 33852 29204
rect 33068 28084 33124 28094
rect 33068 27990 33124 28028
rect 33292 27860 33348 27870
rect 32956 27804 33124 27860
rect 32060 27766 32116 27804
rect 31948 27636 32004 27646
rect 32956 27636 33012 27646
rect 31948 27542 32004 27580
rect 32172 27634 33012 27636
rect 32172 27582 32958 27634
rect 33010 27582 33012 27634
rect 32172 27580 33012 27582
rect 32060 27524 32116 27534
rect 31948 27300 32004 27310
rect 32060 27300 32116 27468
rect 31948 27298 32116 27300
rect 31948 27246 31950 27298
rect 32002 27246 32116 27298
rect 31948 27244 32116 27246
rect 32172 27298 32228 27580
rect 32956 27570 33012 27580
rect 32172 27246 32174 27298
rect 32226 27246 32228 27298
rect 31948 27234 32004 27244
rect 32172 27234 32228 27246
rect 32284 27412 32340 27422
rect 33068 27412 33124 27804
rect 32284 26908 32340 27356
rect 32844 27356 33124 27412
rect 33180 27858 33348 27860
rect 33180 27806 33294 27858
rect 33346 27806 33348 27858
rect 33180 27804 33348 27806
rect 32844 27074 32900 27356
rect 32956 27188 33012 27198
rect 33180 27188 33236 27804
rect 33292 27794 33348 27804
rect 32956 27186 33236 27188
rect 32956 27134 32958 27186
rect 33010 27134 33236 27186
rect 32956 27132 33236 27134
rect 32956 27122 33012 27132
rect 33292 27076 33348 27086
rect 33404 27076 33460 29148
rect 33852 29138 33908 29148
rect 33516 27858 33572 27870
rect 33516 27806 33518 27858
rect 33570 27806 33572 27858
rect 33516 27300 33572 27806
rect 33516 27234 33572 27244
rect 33852 27860 33908 27870
rect 33852 27298 33908 27804
rect 33852 27246 33854 27298
rect 33906 27246 33908 27298
rect 33852 27234 33908 27246
rect 32844 27022 32846 27074
rect 32898 27022 32900 27074
rect 32844 27010 32900 27022
rect 33180 27074 33460 27076
rect 33180 27022 33294 27074
rect 33346 27022 33460 27074
rect 33180 27020 33460 27022
rect 32172 26852 32340 26908
rect 33068 26964 33124 27002
rect 33068 26898 33124 26908
rect 31836 24894 31838 24946
rect 31890 24894 31892 24946
rect 31836 24882 31892 24894
rect 32060 26292 32116 26302
rect 31388 24724 31444 24734
rect 31388 24630 31444 24668
rect 32060 23604 32116 26236
rect 32172 25618 32228 26852
rect 32732 26850 32788 26862
rect 32732 26798 32734 26850
rect 32786 26798 32788 26850
rect 32620 26516 32676 26526
rect 32284 26460 32620 26516
rect 32284 26290 32340 26460
rect 32620 26450 32676 26460
rect 32284 26238 32286 26290
rect 32338 26238 32340 26290
rect 32284 26226 32340 26238
rect 32732 26068 32788 26798
rect 32844 26852 32900 26862
rect 32900 26796 33012 26852
rect 32844 26786 32900 26796
rect 32956 26404 33012 26796
rect 33068 26404 33124 26414
rect 32956 26402 33124 26404
rect 32956 26350 33070 26402
rect 33122 26350 33124 26402
rect 32956 26348 33124 26350
rect 33068 26338 33124 26348
rect 32732 25732 32788 26012
rect 32172 25566 32174 25618
rect 32226 25566 32228 25618
rect 32172 25554 32228 25566
rect 32396 25676 33012 25732
rect 32172 25396 32228 25406
rect 32172 24836 32228 25340
rect 32284 24836 32340 24846
rect 32172 24834 32340 24836
rect 32172 24782 32286 24834
rect 32338 24782 32340 24834
rect 32172 24780 32340 24782
rect 32284 24770 32340 24780
rect 32396 24722 32452 25676
rect 32956 25618 33012 25676
rect 32956 25566 32958 25618
rect 33010 25566 33012 25618
rect 32956 25554 33012 25566
rect 32508 25508 32564 25518
rect 32508 25506 32676 25508
rect 32508 25454 32510 25506
rect 32562 25454 32676 25506
rect 32508 25452 32676 25454
rect 32508 25442 32564 25452
rect 32396 24670 32398 24722
rect 32450 24670 32452 24722
rect 32396 24658 32452 24670
rect 32060 23538 32116 23548
rect 31276 22484 31332 22494
rect 31276 20802 31332 22428
rect 31724 21700 31780 21710
rect 31612 21644 31724 21700
rect 31500 21588 31556 21598
rect 31276 20750 31278 20802
rect 31330 20750 31332 20802
rect 31276 20738 31332 20750
rect 31388 21586 31556 21588
rect 31388 21534 31502 21586
rect 31554 21534 31556 21586
rect 31388 21532 31556 21534
rect 31388 20020 31444 21532
rect 31500 21522 31556 21532
rect 31500 21362 31556 21374
rect 31500 21310 31502 21362
rect 31554 21310 31556 21362
rect 31500 20802 31556 21310
rect 31500 20750 31502 20802
rect 31554 20750 31556 20802
rect 31500 20738 31556 20750
rect 31612 20802 31668 21644
rect 31724 21634 31780 21644
rect 32172 21698 32228 21710
rect 32172 21646 32174 21698
rect 32226 21646 32228 21698
rect 32172 21588 32228 21646
rect 31836 21364 31892 21374
rect 32172 21364 32228 21532
rect 31836 21362 32228 21364
rect 31836 21310 31838 21362
rect 31890 21310 32228 21362
rect 31836 21308 32228 21310
rect 32508 21586 32564 21598
rect 32508 21534 32510 21586
rect 32562 21534 32564 21586
rect 31836 21298 31892 21308
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 31612 20738 31668 20750
rect 31724 20802 31780 20814
rect 31724 20750 31726 20802
rect 31778 20750 31780 20802
rect 31388 19954 31444 19964
rect 31276 19906 31332 19918
rect 31276 19854 31278 19906
rect 31330 19854 31332 19906
rect 31276 19572 31332 19854
rect 31724 19796 31780 20750
rect 31836 20580 31892 20590
rect 31836 20018 31892 20524
rect 31836 19966 31838 20018
rect 31890 19966 31892 20018
rect 31836 19954 31892 19966
rect 31948 19796 32004 21308
rect 32172 20802 32228 20814
rect 32172 20750 32174 20802
rect 32226 20750 32228 20802
rect 32060 20020 32116 20030
rect 32172 20020 32228 20750
rect 32508 20804 32564 21534
rect 32508 20738 32564 20748
rect 32620 20692 32676 25452
rect 32956 25172 33012 25182
rect 32956 24724 33012 25116
rect 33180 24948 33236 27020
rect 33292 27010 33348 27020
rect 33740 26964 33796 26974
rect 33292 26516 33348 26554
rect 33292 26450 33348 26460
rect 33292 26292 33348 26302
rect 33292 26198 33348 26236
rect 33516 26066 33572 26078
rect 33516 26014 33518 26066
rect 33570 26014 33572 26066
rect 33292 25394 33348 25406
rect 33292 25342 33294 25394
rect 33346 25342 33348 25394
rect 33292 25172 33348 25342
rect 33292 25106 33348 25116
rect 33404 24948 33460 24958
rect 33180 24946 33460 24948
rect 33180 24894 33406 24946
rect 33458 24894 33460 24946
rect 33180 24892 33460 24894
rect 33404 24882 33460 24892
rect 33516 24946 33572 26014
rect 33740 25844 33796 26908
rect 33516 24894 33518 24946
rect 33570 24894 33572 24946
rect 33516 24882 33572 24894
rect 33628 25788 33796 25844
rect 33852 26290 33908 26302
rect 33852 26238 33854 26290
rect 33906 26238 33908 26290
rect 33628 24946 33684 25788
rect 33628 24894 33630 24946
rect 33682 24894 33684 24946
rect 33628 24882 33684 24894
rect 33740 25506 33796 25518
rect 33740 25454 33742 25506
rect 33794 25454 33796 25506
rect 32956 24630 33012 24668
rect 33740 23828 33796 25454
rect 33852 25396 33908 26238
rect 34076 25618 34132 29820
rect 34076 25566 34078 25618
rect 34130 25566 34132 25618
rect 34076 25554 34132 25566
rect 33852 25330 33908 25340
rect 33628 23772 33796 23828
rect 34076 24052 34132 24062
rect 33628 22708 33684 23772
rect 33740 23604 33796 23614
rect 33796 23548 33908 23604
rect 33740 23538 33796 23548
rect 32844 22652 33684 22708
rect 33740 23268 33796 23278
rect 32732 22258 32788 22270
rect 32732 22206 32734 22258
rect 32786 22206 32788 22258
rect 32732 21588 32788 22206
rect 32732 21522 32788 21532
rect 32508 20020 32564 20030
rect 32060 20018 32452 20020
rect 32060 19966 32062 20018
rect 32114 19966 32452 20018
rect 32060 19964 32452 19966
rect 32060 19954 32116 19964
rect 32284 19796 32340 19806
rect 31948 19794 32340 19796
rect 31948 19742 32286 19794
rect 32338 19742 32340 19794
rect 31948 19740 32340 19742
rect 31724 19730 31780 19740
rect 32284 19730 32340 19740
rect 31276 19506 31332 19516
rect 31276 19124 31332 19134
rect 31276 19030 31332 19068
rect 31612 19122 31668 19134
rect 31612 19070 31614 19122
rect 31666 19070 31668 19122
rect 31500 17668 31556 17678
rect 31612 17668 31668 19070
rect 31948 19010 32004 19022
rect 31948 18958 31950 19010
rect 32002 18958 32004 19010
rect 31836 17668 31892 17678
rect 31556 17666 31892 17668
rect 31556 17614 31838 17666
rect 31890 17614 31892 17666
rect 31556 17612 31892 17614
rect 31164 17556 31220 17566
rect 31164 17462 31220 17500
rect 31500 17554 31556 17612
rect 31836 17602 31892 17612
rect 31500 17502 31502 17554
rect 31554 17502 31556 17554
rect 31500 17490 31556 17502
rect 31948 16996 32004 18958
rect 32396 17666 32452 19964
rect 32508 19926 32564 19964
rect 32620 19236 32676 20636
rect 32508 19234 32676 19236
rect 32508 19182 32622 19234
rect 32674 19182 32676 19234
rect 32508 19180 32676 19182
rect 32508 18452 32564 19180
rect 32620 19170 32676 19180
rect 32844 18564 32900 22652
rect 33740 22596 33796 23212
rect 33628 22594 33796 22596
rect 33628 22542 33742 22594
rect 33794 22542 33796 22594
rect 33628 22540 33796 22542
rect 33404 22484 33460 22494
rect 33404 22390 33460 22428
rect 33292 22372 33348 22382
rect 33180 22316 33292 22372
rect 33068 22260 33124 22270
rect 33068 22166 33124 22204
rect 33180 22036 33236 22316
rect 33292 22306 33348 22316
rect 33068 21980 33236 22036
rect 33404 22148 33460 22158
rect 33068 21698 33124 21980
rect 33068 21646 33070 21698
rect 33122 21646 33124 21698
rect 33068 21634 33124 21646
rect 33404 21698 33460 22092
rect 33516 22146 33572 22158
rect 33516 22094 33518 22146
rect 33570 22094 33572 22146
rect 33516 22036 33572 22094
rect 33516 21970 33572 21980
rect 33404 21646 33406 21698
rect 33458 21646 33460 21698
rect 33404 21634 33460 21646
rect 33180 21588 33236 21626
rect 33180 21522 33236 21532
rect 33628 21586 33684 22540
rect 33740 22530 33796 22540
rect 33628 21534 33630 21586
rect 33682 21534 33684 21586
rect 33628 21522 33684 21534
rect 33852 21588 33908 23548
rect 34076 22036 34132 23996
rect 34188 23380 34244 31276
rect 34412 31836 34636 31892
rect 34412 30098 34468 31836
rect 34636 31798 34692 31836
rect 34636 30324 34692 30334
rect 34748 30324 34804 32398
rect 35308 32452 35364 32462
rect 35644 32452 35700 32462
rect 35308 32450 35588 32452
rect 35308 32398 35310 32450
rect 35362 32398 35588 32450
rect 35308 32396 35588 32398
rect 35308 32386 35364 32396
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35308 31666 35364 31678
rect 35308 31614 35310 31666
rect 35362 31614 35364 31666
rect 35308 31556 35364 31614
rect 35308 31490 35364 31500
rect 35532 31218 35588 32396
rect 35644 32358 35700 32396
rect 35756 31780 35812 31790
rect 35756 31686 35812 31724
rect 35980 31780 36036 32510
rect 35980 31714 36036 31724
rect 36204 31778 36260 31790
rect 36204 31726 36206 31778
rect 36258 31726 36260 31778
rect 35532 31166 35534 31218
rect 35586 31166 35588 31218
rect 35532 31154 35588 31166
rect 35868 31220 35924 31230
rect 35868 31126 35924 31164
rect 35084 31108 35140 31118
rect 35308 31108 35364 31118
rect 35140 31106 35364 31108
rect 35140 31054 35310 31106
rect 35362 31054 35364 31106
rect 35140 31052 35364 31054
rect 35084 31014 35140 31052
rect 35308 31042 35364 31052
rect 35756 30996 35812 31006
rect 35756 30994 35924 30996
rect 35756 30942 35758 30994
rect 35810 30942 35924 30994
rect 35756 30940 35924 30942
rect 35756 30930 35812 30940
rect 35644 30884 35700 30894
rect 35644 30790 35700 30828
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34692 30268 34804 30324
rect 35868 30324 35924 30940
rect 34636 30230 34692 30268
rect 34412 30046 34414 30098
rect 34466 30046 34468 30098
rect 34412 28420 34468 30046
rect 34524 30100 34580 30110
rect 34524 30006 34580 30044
rect 35532 29426 35588 29438
rect 35532 29374 35534 29426
rect 35586 29374 35588 29426
rect 35532 29204 35588 29374
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35420 28644 35476 28654
rect 35532 28644 35588 29148
rect 35420 28642 35588 28644
rect 35420 28590 35422 28642
rect 35474 28590 35588 28642
rect 35420 28588 35588 28590
rect 35644 29428 35700 29438
rect 35420 28578 35476 28588
rect 34412 28354 34468 28364
rect 35532 28420 35588 28430
rect 35532 28326 35588 28364
rect 35420 27746 35476 27758
rect 35420 27694 35422 27746
rect 35474 27694 35476 27746
rect 35420 27636 35476 27694
rect 35420 27570 35476 27580
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35308 27300 35364 27310
rect 35308 27206 35364 27244
rect 34860 27188 34916 27198
rect 34860 27094 34916 27132
rect 34300 27076 34356 27086
rect 34748 27076 34804 27086
rect 34300 27074 34468 27076
rect 34300 27022 34302 27074
rect 34354 27022 34468 27074
rect 34300 27020 34468 27022
rect 34300 27010 34356 27020
rect 34412 25620 34468 27020
rect 34524 26964 34580 27002
rect 34524 26898 34580 26908
rect 34748 26962 34804 27020
rect 35420 27076 35476 27086
rect 35420 26982 35476 27020
rect 34748 26910 34750 26962
rect 34802 26910 34804 26962
rect 34748 26908 34804 26910
rect 34748 26852 34916 26908
rect 34860 26402 34916 26852
rect 34860 26350 34862 26402
rect 34914 26350 34916 26402
rect 34860 26338 34916 26350
rect 35308 26180 35364 26190
rect 35308 26086 35364 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34748 25620 34804 25630
rect 34412 25618 34804 25620
rect 34412 25566 34750 25618
rect 34802 25566 34804 25618
rect 34412 25564 34804 25566
rect 34748 25554 34804 25564
rect 35644 25618 35700 29372
rect 35868 29428 35924 30268
rect 36204 30324 36260 31726
rect 36316 31556 36372 32844
rect 36428 32004 36484 33292
rect 36540 33124 36596 33134
rect 37100 33124 37156 33134
rect 37772 33124 37828 33134
rect 36540 33122 37044 33124
rect 36540 33070 36542 33122
rect 36594 33070 37044 33122
rect 36540 33068 37044 33070
rect 36540 33058 36596 33068
rect 36988 32788 37044 33068
rect 37100 33122 37268 33124
rect 37100 33070 37102 33122
rect 37154 33070 37268 33122
rect 37100 33068 37268 33070
rect 37100 33058 37156 33068
rect 37100 32788 37156 32798
rect 36988 32786 37156 32788
rect 36988 32734 37102 32786
rect 37154 32734 37156 32786
rect 36988 32732 37156 32734
rect 37100 32722 37156 32732
rect 36652 32564 36708 32574
rect 36652 32470 36708 32508
rect 36876 32562 36932 32574
rect 36876 32510 36878 32562
rect 36930 32510 36932 32562
rect 36876 32228 36932 32510
rect 37100 32564 37156 32574
rect 37212 32564 37268 33068
rect 37772 32674 37828 33068
rect 37772 32622 37774 32674
rect 37826 32622 37828 32674
rect 37772 32610 37828 32622
rect 37156 32508 37268 32564
rect 37324 32564 37380 32574
rect 37660 32564 37716 32574
rect 37324 32562 37716 32564
rect 37324 32510 37326 32562
rect 37378 32510 37662 32562
rect 37714 32510 37716 32562
rect 37324 32508 37716 32510
rect 37100 32498 37156 32508
rect 37324 32498 37380 32508
rect 37660 32498 37716 32508
rect 36428 31938 36484 31948
rect 36764 32172 36932 32228
rect 36988 32450 37044 32462
rect 36988 32398 36990 32450
rect 37042 32398 37044 32450
rect 36764 31892 36820 32172
rect 36316 31490 36372 31500
rect 36540 31668 36596 31678
rect 36316 31332 36372 31342
rect 36316 30994 36372 31276
rect 36540 31218 36596 31612
rect 36540 31166 36542 31218
rect 36594 31166 36596 31218
rect 36540 31154 36596 31166
rect 36316 30942 36318 30994
rect 36370 30942 36372 30994
rect 36316 30930 36372 30942
rect 36652 30770 36708 30782
rect 36652 30718 36654 30770
rect 36706 30718 36708 30770
rect 36316 30324 36372 30334
rect 36204 30322 36372 30324
rect 36204 30270 36318 30322
rect 36370 30270 36372 30322
rect 36204 30268 36372 30270
rect 36204 30212 36260 30268
rect 36316 30258 36372 30268
rect 35980 29988 36036 29998
rect 35980 29894 36036 29932
rect 36092 29652 36148 29662
rect 36204 29652 36260 30156
rect 36092 29650 36260 29652
rect 36092 29598 36094 29650
rect 36146 29598 36260 29650
rect 36092 29596 36260 29598
rect 36428 29988 36484 29998
rect 36652 29988 36708 30718
rect 36764 30548 36820 31836
rect 36876 32004 36932 32014
rect 36876 31778 36932 31948
rect 36988 31892 37044 32398
rect 36988 31826 37044 31836
rect 37884 31892 37940 31902
rect 37884 31798 37940 31836
rect 36876 31726 36878 31778
rect 36930 31726 36932 31778
rect 36876 31714 36932 31726
rect 37100 31780 37156 31790
rect 37100 31686 37156 31724
rect 37212 31778 37268 31790
rect 37212 31726 37214 31778
rect 37266 31726 37268 31778
rect 37212 31556 37268 31726
rect 38220 31778 38276 31790
rect 38220 31726 38222 31778
rect 38274 31726 38276 31778
rect 37548 31668 37604 31678
rect 37548 31574 37604 31612
rect 37212 31490 37268 31500
rect 37996 31554 38052 31566
rect 37996 31502 37998 31554
rect 38050 31502 38052 31554
rect 37996 31106 38052 31502
rect 38220 31556 38276 31726
rect 38668 31556 38724 31566
rect 38220 31554 38724 31556
rect 38220 31502 38670 31554
rect 38722 31502 38724 31554
rect 38220 31500 38724 31502
rect 37996 31054 37998 31106
rect 38050 31054 38052 31106
rect 37996 31042 38052 31054
rect 37212 30994 37268 31006
rect 37212 30942 37214 30994
rect 37266 30942 37268 30994
rect 36764 30492 37044 30548
rect 36988 30098 37044 30492
rect 36988 30046 36990 30098
rect 37042 30046 37044 30098
rect 36988 30034 37044 30046
rect 36428 29986 36708 29988
rect 36428 29934 36430 29986
rect 36482 29934 36708 29986
rect 36428 29932 36708 29934
rect 36876 29988 36932 29998
rect 36092 29586 36148 29596
rect 35868 29334 35924 29372
rect 35980 29314 36036 29326
rect 35980 29262 35982 29314
rect 36034 29262 36036 29314
rect 35756 28418 35812 28430
rect 35756 28366 35758 28418
rect 35810 28366 35812 28418
rect 35756 27860 35812 28366
rect 35868 27860 35924 27870
rect 35756 27858 35924 27860
rect 35756 27806 35870 27858
rect 35922 27806 35924 27858
rect 35756 27804 35924 27806
rect 35868 27794 35924 27804
rect 35980 27074 36036 29262
rect 36316 27746 36372 27758
rect 36316 27694 36318 27746
rect 36370 27694 36372 27746
rect 36316 27300 36372 27694
rect 36316 27234 36372 27244
rect 35980 27022 35982 27074
rect 36034 27022 36036 27074
rect 35980 27010 36036 27022
rect 36316 26852 36372 26862
rect 36316 26402 36372 26796
rect 36316 26350 36318 26402
rect 36370 26350 36372 26402
rect 36316 26338 36372 26350
rect 35644 25566 35646 25618
rect 35698 25566 35700 25618
rect 35644 25554 35700 25566
rect 35756 26290 35812 26302
rect 35756 26238 35758 26290
rect 35810 26238 35812 26290
rect 35196 25508 35252 25518
rect 34188 23314 34244 23324
rect 35084 25506 35252 25508
rect 35084 25454 35198 25506
rect 35250 25454 35252 25506
rect 35084 25452 35252 25454
rect 34412 23266 34468 23278
rect 34412 23214 34414 23266
rect 34466 23214 34468 23266
rect 34300 23156 34356 23166
rect 34188 23154 34356 23156
rect 34188 23102 34302 23154
rect 34354 23102 34356 23154
rect 34188 23100 34356 23102
rect 34188 22372 34244 23100
rect 34300 23090 34356 23100
rect 34188 22258 34244 22316
rect 34188 22206 34190 22258
rect 34242 22206 34244 22258
rect 34188 22194 34244 22206
rect 34412 22260 34468 23214
rect 34636 23156 34692 23166
rect 34636 23154 35028 23156
rect 34636 23102 34638 23154
rect 34690 23102 35028 23154
rect 34636 23100 35028 23102
rect 34636 23090 34692 23100
rect 34412 22166 34468 22204
rect 34524 22146 34580 22158
rect 34524 22094 34526 22146
rect 34578 22094 34580 22146
rect 34076 21980 34356 22036
rect 33852 21522 33908 21532
rect 33292 21476 33348 21486
rect 33292 20690 33348 21420
rect 34188 21476 34244 21486
rect 34188 21382 34244 21420
rect 33292 20638 33294 20690
rect 33346 20638 33348 20690
rect 33292 20580 33348 20638
rect 33852 21362 33908 21374
rect 33852 21310 33854 21362
rect 33906 21310 33908 21362
rect 33292 20514 33348 20524
rect 33628 20578 33684 20590
rect 33628 20526 33630 20578
rect 33682 20526 33684 20578
rect 33404 20242 33460 20254
rect 33404 20190 33406 20242
rect 33458 20190 33460 20242
rect 33404 20132 33460 20190
rect 33404 20066 33460 20076
rect 32956 20020 33012 20030
rect 32956 19124 33012 19964
rect 33516 20020 33572 20030
rect 33516 19926 33572 19964
rect 32956 19030 33012 19068
rect 33628 18900 33684 20526
rect 33852 20356 33908 21310
rect 34188 20804 34244 20814
rect 34300 20804 34356 21980
rect 34244 20748 34356 20804
rect 34188 20710 34244 20748
rect 34524 20580 34580 22094
rect 34636 22148 34692 22158
rect 34636 22054 34692 22092
rect 34860 21700 34916 21710
rect 34860 21606 34916 21644
rect 34748 20692 34804 20702
rect 34748 20598 34804 20636
rect 34524 20514 34580 20524
rect 33852 20290 33908 20300
rect 34188 20356 34244 20366
rect 33740 20020 33796 20030
rect 33740 19926 33796 19964
rect 34076 20018 34132 20030
rect 34076 19966 34078 20018
rect 34130 19966 34132 20018
rect 33852 19796 33908 19806
rect 34076 19796 34132 19966
rect 33628 18834 33684 18844
rect 33740 19740 33852 19796
rect 33908 19740 34132 19796
rect 34188 19908 34244 20300
rect 34748 20244 34804 20254
rect 34412 20242 34804 20244
rect 34412 20190 34750 20242
rect 34802 20190 34804 20242
rect 34412 20188 34804 20190
rect 34300 20132 34356 20142
rect 34412 20132 34468 20188
rect 34748 20178 34804 20188
rect 34300 20130 34468 20132
rect 34300 20078 34302 20130
rect 34354 20078 34468 20130
rect 34300 20076 34468 20078
rect 34300 20066 34356 20076
rect 34636 20074 34692 20086
rect 34636 20022 34638 20074
rect 34690 20022 34692 20074
rect 34636 19908 34692 20022
rect 34188 19852 34692 19908
rect 34860 20020 34916 20030
rect 34972 20020 35028 23100
rect 35084 21700 35140 25452
rect 35196 25442 35252 25452
rect 35756 24612 35812 26238
rect 36428 26290 36484 29932
rect 36876 29428 36932 29932
rect 37212 29428 37268 30942
rect 37660 30884 37716 30894
rect 37660 30434 37716 30828
rect 37660 30382 37662 30434
rect 37714 30382 37716 30434
rect 37660 30370 37716 30382
rect 37996 30322 38052 30334
rect 37996 30270 37998 30322
rect 38050 30270 38052 30322
rect 37324 30212 37380 30222
rect 37324 30118 37380 30156
rect 37884 29988 37940 29998
rect 37884 29540 37940 29932
rect 37884 29474 37940 29484
rect 37996 29538 38052 30270
rect 38444 29988 38500 31500
rect 38668 31490 38724 31500
rect 40124 30882 40180 30894
rect 40124 30830 40126 30882
rect 40178 30830 40180 30882
rect 40124 30324 40180 30830
rect 40124 30258 40180 30268
rect 38444 29894 38500 29932
rect 37996 29486 37998 29538
rect 38050 29486 38052 29538
rect 37996 29474 38052 29486
rect 36876 29426 37268 29428
rect 36876 29374 37214 29426
rect 37266 29374 37268 29426
rect 36876 29372 37268 29374
rect 36876 29314 36932 29372
rect 37212 29362 37268 29372
rect 38220 29428 38276 29438
rect 36876 29262 36878 29314
rect 36930 29262 36932 29314
rect 36428 26238 36430 26290
rect 36482 26238 36484 26290
rect 36428 26226 36484 26238
rect 36764 26290 36820 26302
rect 36764 26238 36766 26290
rect 36818 26238 36820 26290
rect 35644 24556 35756 24612
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35644 22596 35700 24556
rect 35756 24546 35812 24556
rect 36764 24052 36820 26238
rect 36876 24948 36932 29262
rect 38220 28530 38276 29372
rect 38220 28478 38222 28530
rect 38274 28478 38276 28530
rect 38220 28466 38276 28478
rect 38556 29316 38612 29326
rect 38556 28642 38612 29260
rect 40124 29316 40180 29326
rect 40124 29222 40180 29260
rect 38556 28590 38558 28642
rect 38610 28590 38612 28642
rect 37996 27300 38052 27310
rect 37996 27206 38052 27244
rect 38556 27186 38612 28590
rect 38556 27134 38558 27186
rect 38610 27134 38612 27186
rect 38556 27122 38612 27134
rect 38332 27074 38388 27086
rect 38332 27022 38334 27074
rect 38386 27022 38388 27074
rect 36876 24946 37268 24948
rect 36876 24894 36878 24946
rect 36930 24894 37268 24946
rect 36876 24892 37268 24894
rect 36876 24882 36932 24892
rect 36764 23986 36820 23996
rect 37212 24722 37268 24892
rect 37212 24670 37214 24722
rect 37266 24670 37268 24722
rect 36540 23940 36596 23950
rect 36540 23846 36596 23884
rect 37212 23940 37268 24670
rect 37996 24612 38052 24622
rect 37212 23846 37268 23884
rect 37548 24610 38052 24612
rect 37548 24558 37998 24610
rect 38050 24558 38052 24610
rect 37548 24556 38052 24558
rect 36652 23380 36708 23390
rect 36652 23286 36708 23324
rect 37548 23378 37604 24556
rect 37996 24546 38052 24556
rect 37996 23828 38052 23838
rect 37548 23326 37550 23378
rect 37602 23326 37604 23378
rect 37548 23314 37604 23326
rect 37660 23826 38052 23828
rect 37660 23774 37998 23826
rect 38050 23774 38052 23826
rect 37660 23772 38052 23774
rect 35308 22540 35700 22596
rect 36316 23266 36372 23278
rect 36316 23214 36318 23266
rect 36370 23214 36372 23266
rect 35308 22372 35364 22540
rect 35084 21634 35140 21644
rect 35196 22370 35364 22372
rect 35196 22318 35310 22370
rect 35362 22318 35364 22370
rect 35196 22316 35364 22318
rect 35196 22036 35252 22316
rect 35308 22306 35364 22316
rect 35532 22372 35588 22382
rect 35532 22258 35588 22316
rect 35532 22206 35534 22258
rect 35586 22206 35588 22258
rect 35532 22194 35588 22206
rect 35868 22370 35924 22382
rect 35868 22318 35870 22370
rect 35922 22318 35924 22370
rect 35868 22260 35924 22318
rect 35196 21698 35252 21980
rect 35196 21646 35198 21698
rect 35250 21646 35252 21698
rect 35196 21634 35252 21646
rect 35532 21700 35588 21710
rect 35420 21588 35476 21598
rect 35420 21494 35476 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20020 35140 20030
rect 34972 20018 35140 20020
rect 34972 19966 35086 20018
rect 35138 19966 35140 20018
rect 34972 19964 35140 19966
rect 32508 18386 32564 18396
rect 32620 18508 32900 18564
rect 33740 18674 33796 19740
rect 33852 19730 33908 19740
rect 33740 18622 33742 18674
rect 33794 18622 33796 18674
rect 33740 18564 33796 18622
rect 32396 17614 32398 17666
rect 32450 17614 32452 17666
rect 32396 17602 32452 17614
rect 32620 17556 32676 18508
rect 33740 18498 33796 18508
rect 34076 18450 34132 18462
rect 34076 18398 34078 18450
rect 34130 18398 34132 18450
rect 34076 18228 34132 18398
rect 34076 18162 34132 18172
rect 34188 17780 34244 19852
rect 34412 19124 34468 19134
rect 33964 17724 34244 17780
rect 34300 18452 34356 18462
rect 33964 17666 34020 17724
rect 33964 17614 33966 17666
rect 34018 17614 34020 17666
rect 32508 17554 32676 17556
rect 32508 17502 32622 17554
rect 32674 17502 32676 17554
rect 32508 17500 32676 17502
rect 32172 17444 32228 17454
rect 32172 17350 32228 17388
rect 31948 16930 32004 16940
rect 32508 16772 32564 17500
rect 32620 17490 32676 17500
rect 32732 17556 32788 17566
rect 33068 17556 33124 17566
rect 32732 17554 33012 17556
rect 32732 17502 32734 17554
rect 32786 17502 33012 17554
rect 32732 17500 33012 17502
rect 32732 17490 32788 17500
rect 31612 16716 32564 16772
rect 32844 16772 32900 16782
rect 31612 16098 31668 16716
rect 31612 16046 31614 16098
rect 31666 16046 31668 16098
rect 31612 16034 31668 16046
rect 31948 15988 32004 15998
rect 31724 15932 31948 15988
rect 31276 15484 31556 15540
rect 31052 15250 31108 15260
rect 31164 15314 31220 15326
rect 31164 15262 31166 15314
rect 31218 15262 31220 15314
rect 31052 15092 31108 15102
rect 31052 14998 31108 15036
rect 31164 14980 31220 15262
rect 31164 14914 31220 14924
rect 30940 14802 30996 14812
rect 30828 14642 31220 14644
rect 30828 14590 30830 14642
rect 30882 14590 31220 14642
rect 30828 14588 31220 14590
rect 30828 14578 30884 14588
rect 31164 14530 31220 14588
rect 31164 14478 31166 14530
rect 31218 14478 31220 14530
rect 31164 14466 31220 14478
rect 30716 13972 30772 13982
rect 30604 13970 30772 13972
rect 30604 13918 30718 13970
rect 30770 13918 30772 13970
rect 30604 13916 30772 13918
rect 30716 13906 30772 13916
rect 31164 13748 31220 13758
rect 31276 13748 31332 15484
rect 31500 15428 31556 15484
rect 31612 15428 31668 15438
rect 31724 15428 31780 15932
rect 31948 15894 32004 15932
rect 31500 15426 31780 15428
rect 31500 15374 31614 15426
rect 31666 15374 31780 15426
rect 31500 15372 31780 15374
rect 31612 15362 31668 15372
rect 30492 13692 30884 13748
rect 30716 13524 30772 13534
rect 30268 13468 30660 13524
rect 30268 12850 30324 13468
rect 30604 13412 30660 13468
rect 30604 13346 30660 13356
rect 30716 12962 30772 13468
rect 30716 12910 30718 12962
rect 30770 12910 30772 12962
rect 30716 12898 30772 12910
rect 30828 13300 30884 13692
rect 31164 13746 31332 13748
rect 31164 13694 31166 13746
rect 31218 13694 31332 13746
rect 31164 13692 31332 13694
rect 31388 15316 31444 15326
rect 31388 13746 31444 15260
rect 31388 13694 31390 13746
rect 31442 13694 31444 13746
rect 31164 13682 31220 13692
rect 31388 13412 31444 13694
rect 31612 14980 31668 14990
rect 31612 13860 31668 14924
rect 32060 14756 32116 16716
rect 32844 15540 32900 16716
rect 32844 15474 32900 15484
rect 32956 15428 33012 17500
rect 33068 16994 33124 17500
rect 33852 17556 33908 17566
rect 33852 17462 33908 17500
rect 33404 17108 33460 17118
rect 33852 17108 33908 17118
rect 33404 17014 33460 17052
rect 33740 17052 33852 17108
rect 33964 17108 34020 17614
rect 34076 17556 34132 17566
rect 34076 17554 34244 17556
rect 34076 17502 34078 17554
rect 34130 17502 34244 17554
rect 34076 17500 34244 17502
rect 34076 17490 34132 17500
rect 34076 17108 34132 17118
rect 33964 17106 34132 17108
rect 33964 17054 34078 17106
rect 34130 17054 34132 17106
rect 33964 17052 34132 17054
rect 33068 16942 33070 16994
rect 33122 16942 33124 16994
rect 33068 15988 33124 16942
rect 33516 16772 33572 16782
rect 33516 16324 33572 16716
rect 33068 15922 33124 15932
rect 33404 16322 33572 16324
rect 33404 16270 33518 16322
rect 33570 16270 33572 16322
rect 33404 16268 33572 16270
rect 33180 15874 33236 15886
rect 33180 15822 33182 15874
rect 33234 15822 33236 15874
rect 33180 15652 33236 15822
rect 33292 15652 33348 15662
rect 33180 15596 33292 15652
rect 33068 15428 33124 15438
rect 32956 15426 33124 15428
rect 32956 15374 33070 15426
rect 33122 15374 33124 15426
rect 32956 15372 33124 15374
rect 32172 15316 32228 15326
rect 32172 15222 32228 15260
rect 32060 14690 32116 14700
rect 32172 15090 32228 15102
rect 32508 15092 32564 15102
rect 32172 15038 32174 15090
rect 32226 15038 32228 15090
rect 32172 14084 32228 15038
rect 32172 14018 32228 14028
rect 32284 15090 32564 15092
rect 32284 15038 32510 15090
rect 32562 15038 32564 15090
rect 32284 15036 32564 15038
rect 32172 13860 32228 13870
rect 31612 13858 32228 13860
rect 31612 13806 32174 13858
rect 32226 13806 32228 13858
rect 31612 13804 32228 13806
rect 31612 13746 31668 13804
rect 31612 13694 31614 13746
rect 31666 13694 31668 13746
rect 31612 13524 31668 13694
rect 31612 13458 31668 13468
rect 31836 13634 31892 13646
rect 31836 13582 31838 13634
rect 31890 13582 31892 13634
rect 31388 13346 31444 13356
rect 30828 13244 31220 13300
rect 30828 12962 30884 13244
rect 31164 13188 31220 13244
rect 31836 13188 31892 13582
rect 31164 13132 31892 13188
rect 30828 12910 30830 12962
rect 30882 12910 30884 12962
rect 30828 12898 30884 12910
rect 31052 12964 31108 12974
rect 31052 12870 31108 12908
rect 31276 12962 31332 12974
rect 31276 12910 31278 12962
rect 31330 12910 31332 12962
rect 30268 12798 30270 12850
rect 30322 12798 30324 12850
rect 30268 12786 30324 12798
rect 31164 12852 31220 12862
rect 30156 12572 30884 12628
rect 29820 12114 29876 12124
rect 29932 12460 30100 12516
rect 27916 11956 27972 11966
rect 28700 11956 28756 11966
rect 27916 11954 28196 11956
rect 27916 11902 27918 11954
rect 27970 11902 28196 11954
rect 27916 11900 28196 11902
rect 27916 11890 27972 11900
rect 28140 11282 28196 11900
rect 28700 11954 29204 11956
rect 28700 11902 28702 11954
rect 28754 11902 29204 11954
rect 28700 11900 29204 11902
rect 28700 11890 28756 11900
rect 29148 11394 29204 11900
rect 29148 11342 29150 11394
rect 29202 11342 29204 11394
rect 28140 11230 28142 11282
rect 28194 11230 28196 11282
rect 28140 11218 28196 11230
rect 28252 11284 28308 11294
rect 28252 11190 28308 11228
rect 27916 11172 27972 11182
rect 27916 11078 27972 11116
rect 28588 11172 28644 11182
rect 27580 10782 27582 10834
rect 27634 10782 27636 10834
rect 27580 10770 27636 10782
rect 28252 10724 28308 10734
rect 27916 10610 27972 10622
rect 27916 10558 27918 10610
rect 27970 10558 27972 10610
rect 27804 9826 27860 9838
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27692 9156 27748 9166
rect 27692 9042 27748 9100
rect 27804 9154 27860 9774
rect 27916 9602 27972 10558
rect 27916 9550 27918 9602
rect 27970 9550 27972 9602
rect 27916 9538 27972 9550
rect 28140 9268 28196 9278
rect 28140 9174 28196 9212
rect 28252 9266 28308 10668
rect 28588 10610 28644 11116
rect 28924 10724 28980 10734
rect 28924 10630 28980 10668
rect 28588 10558 28590 10610
rect 28642 10558 28644 10610
rect 28588 10546 28644 10558
rect 29148 10050 29204 11342
rect 29484 11284 29540 11294
rect 29484 11190 29540 11228
rect 29260 11172 29316 11182
rect 29260 11170 29428 11172
rect 29260 11118 29262 11170
rect 29314 11118 29428 11170
rect 29260 11116 29428 11118
rect 29260 11106 29316 11116
rect 29148 9998 29150 10050
rect 29202 9998 29204 10050
rect 29148 9986 29204 9998
rect 29372 9714 29428 11116
rect 29932 10834 29988 12460
rect 30828 12178 30884 12572
rect 30828 12126 30830 12178
rect 30882 12126 30884 12178
rect 29932 10782 29934 10834
rect 29986 10782 29988 10834
rect 29932 10770 29988 10782
rect 30044 11284 30100 11294
rect 29708 10724 29764 10734
rect 29484 10612 29540 10622
rect 29484 10050 29540 10556
rect 29708 10610 29764 10668
rect 29708 10558 29710 10610
rect 29762 10558 29764 10610
rect 29708 10546 29764 10558
rect 30044 10610 30100 11228
rect 30828 11172 30884 12126
rect 30940 12290 30996 12302
rect 31164 12292 31220 12796
rect 31276 12628 31332 12910
rect 31500 12962 31556 13132
rect 31948 13076 32004 13804
rect 32172 13794 32228 13804
rect 31500 12910 31502 12962
rect 31554 12910 31556 12962
rect 31500 12898 31556 12910
rect 31836 13020 32004 13076
rect 32060 13636 32116 13646
rect 31836 12962 31892 13020
rect 31836 12910 31838 12962
rect 31890 12910 31892 12962
rect 31836 12898 31892 12910
rect 31724 12850 31780 12862
rect 31724 12798 31726 12850
rect 31778 12798 31780 12850
rect 31724 12628 31780 12798
rect 32060 12628 32116 13580
rect 31276 12572 31780 12628
rect 30940 12238 30942 12290
rect 30994 12238 30996 12290
rect 30940 11396 30996 12238
rect 30940 11330 30996 11340
rect 31052 12290 31220 12292
rect 31052 12238 31166 12290
rect 31218 12238 31220 12290
rect 31052 12236 31220 12238
rect 30828 11106 30884 11116
rect 30044 10558 30046 10610
rect 30098 10558 30100 10610
rect 30044 10546 30100 10558
rect 30268 10612 30324 10622
rect 30268 10518 30324 10556
rect 29484 9998 29486 10050
rect 29538 9998 29540 10050
rect 29484 9986 29540 9998
rect 29372 9662 29374 9714
rect 29426 9662 29428 9714
rect 28252 9214 28254 9266
rect 28306 9214 28308 9266
rect 28252 9202 28308 9214
rect 29148 9268 29204 9278
rect 29148 9174 29204 9212
rect 28588 9156 28644 9166
rect 27804 9102 27806 9154
rect 27858 9102 27860 9154
rect 27804 9090 27860 9102
rect 28476 9154 28644 9156
rect 28476 9102 28590 9154
rect 28642 9102 28644 9154
rect 28476 9100 28644 9102
rect 27692 8990 27694 9042
rect 27746 8990 27748 9042
rect 27692 8978 27748 8990
rect 28364 9042 28420 9054
rect 28364 8990 28366 9042
rect 28418 8990 28420 9042
rect 28364 8708 28420 8990
rect 26460 6690 26516 6748
rect 26460 6638 26462 6690
rect 26514 6638 26516 6690
rect 26460 6626 26516 6638
rect 27132 8372 27300 8428
rect 27804 8652 28420 8708
rect 27132 6468 27188 8372
rect 27804 8370 27860 8652
rect 27804 8318 27806 8370
rect 27858 8318 27860 8370
rect 27804 8306 27860 8318
rect 28252 8484 28308 8494
rect 27580 8258 27636 8270
rect 27580 8206 27582 8258
rect 27634 8206 27636 8258
rect 27580 8036 27636 8206
rect 27916 8260 27972 8270
rect 28252 8260 28308 8428
rect 28364 8484 28420 8494
rect 28476 8484 28532 9100
rect 28588 9090 28644 9100
rect 28364 8482 28532 8484
rect 28364 8430 28366 8482
rect 28418 8430 28532 8482
rect 28364 8428 28532 8430
rect 28364 8418 28420 8428
rect 27916 8258 28308 8260
rect 27916 8206 27918 8258
rect 27970 8206 28254 8258
rect 28306 8206 28308 8258
rect 27916 8204 28308 8206
rect 27916 8194 27972 8204
rect 28252 8194 28308 8204
rect 27580 7970 27636 7980
rect 28364 8036 28420 8046
rect 28364 7942 28420 7980
rect 27468 6916 27524 6926
rect 27468 6690 27524 6860
rect 27468 6638 27470 6690
rect 27522 6638 27524 6690
rect 27468 6626 27524 6638
rect 28364 6916 28420 6926
rect 27132 6374 27188 6412
rect 26348 6290 26404 6300
rect 26236 5966 26238 6018
rect 26290 5966 26292 6018
rect 26236 5954 26292 5966
rect 28364 5794 28420 6860
rect 29372 6916 29428 9662
rect 30940 9940 30996 9950
rect 31052 9940 31108 12236
rect 31164 12226 31220 12236
rect 31612 12180 31668 12190
rect 31612 12086 31668 12124
rect 31724 11284 31780 12572
rect 31836 12572 32116 12628
rect 32172 13188 32228 13198
rect 31836 12402 31892 12572
rect 31836 12350 31838 12402
rect 31890 12350 31892 12402
rect 31836 12338 31892 12350
rect 32172 12404 32228 13132
rect 32284 13188 32340 15036
rect 32508 15026 32564 15036
rect 33068 13860 33124 15372
rect 33068 13794 33124 13804
rect 32508 13746 32564 13758
rect 32508 13694 32510 13746
rect 32562 13694 32564 13746
rect 32508 13636 32564 13694
rect 33180 13636 33236 13646
rect 32508 13634 33236 13636
rect 32508 13582 33182 13634
rect 33234 13582 33236 13634
rect 32508 13580 33236 13582
rect 32508 13412 32564 13580
rect 32508 13346 32564 13356
rect 32844 13188 32900 13198
rect 32284 13186 32900 13188
rect 32284 13134 32286 13186
rect 32338 13134 32846 13186
rect 32898 13134 32900 13186
rect 32284 13132 32900 13134
rect 32284 13122 32340 13132
rect 32844 13122 32900 13132
rect 33068 13188 33124 13198
rect 33068 13094 33124 13132
rect 32620 12964 32676 12974
rect 32620 12870 32676 12908
rect 32732 12738 32788 12750
rect 32732 12686 32734 12738
rect 32786 12686 32788 12738
rect 32284 12404 32340 12414
rect 32172 12402 32340 12404
rect 32172 12350 32286 12402
rect 32338 12350 32340 12402
rect 32172 12348 32340 12350
rect 32284 12338 32340 12348
rect 31724 11218 31780 11228
rect 30940 9938 31108 9940
rect 30940 9886 30942 9938
rect 30994 9886 31108 9938
rect 30940 9884 31108 9886
rect 31388 11172 31444 11182
rect 31388 9938 31444 11116
rect 31836 11172 31892 11182
rect 31948 11172 32004 11182
rect 31892 11170 32004 11172
rect 31892 11118 31950 11170
rect 32002 11118 32004 11170
rect 31892 11116 32004 11118
rect 31836 11106 31892 11116
rect 31948 11106 32004 11116
rect 31388 9886 31390 9938
rect 31442 9886 31444 9938
rect 29596 9604 29652 9614
rect 29596 8930 29652 9548
rect 30380 9604 30436 9614
rect 30380 9510 30436 9548
rect 30940 9268 30996 9884
rect 31388 9828 31444 9886
rect 31388 9762 31444 9772
rect 31724 10388 31780 10398
rect 30940 9202 30996 9212
rect 31724 9154 31780 10332
rect 32732 10388 32788 12686
rect 33180 12402 33236 13580
rect 33292 13188 33348 15596
rect 33404 15538 33460 16268
rect 33516 16258 33572 16268
rect 33740 15986 33796 17052
rect 33852 17042 33908 17052
rect 34076 17042 34132 17052
rect 34188 16772 34244 17500
rect 34300 17332 34356 18396
rect 34412 18450 34468 19068
rect 34636 18564 34692 18574
rect 34860 18564 34916 19964
rect 35084 19954 35140 19964
rect 35420 20020 35476 20030
rect 35420 19926 35476 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34860 18508 35028 18564
rect 34636 18470 34692 18508
rect 34412 18398 34414 18450
rect 34466 18398 34468 18450
rect 34412 18386 34468 18398
rect 34860 18340 34916 18350
rect 34860 18246 34916 18284
rect 34636 18228 34692 18238
rect 34524 17892 34580 17902
rect 34524 17798 34580 17836
rect 34300 16772 34356 17276
rect 34636 16996 34692 18172
rect 34636 16882 34692 16940
rect 34972 17108 35028 18508
rect 35084 18450 35140 18462
rect 35084 18398 35086 18450
rect 35138 18398 35140 18450
rect 35084 17780 35140 18398
rect 35308 18338 35364 18350
rect 35308 18286 35310 18338
rect 35362 18286 35364 18338
rect 35308 18228 35364 18286
rect 35532 18340 35588 21644
rect 35868 21586 35924 22204
rect 36204 22258 36260 22270
rect 36204 22206 36206 22258
rect 36258 22206 36260 22258
rect 36092 22146 36148 22158
rect 36092 22094 36094 22146
rect 36146 22094 36148 22146
rect 36092 21700 36148 22094
rect 36092 21634 36148 21644
rect 35868 21534 35870 21586
rect 35922 21534 35924 21586
rect 35868 21522 35924 21534
rect 36092 21364 36148 21374
rect 36204 21364 36260 22206
rect 36316 22148 36372 23214
rect 37436 23266 37492 23278
rect 37436 23214 37438 23266
rect 37490 23214 37492 23266
rect 37324 22372 37380 22382
rect 37324 22278 37380 22316
rect 36316 22082 36372 22092
rect 36876 22148 36932 22158
rect 36428 21812 36484 21822
rect 36428 21718 36484 21756
rect 36092 21362 36260 21364
rect 36092 21310 36094 21362
rect 36146 21310 36260 21362
rect 36092 21308 36260 21310
rect 36092 18450 36148 21308
rect 36428 20578 36484 20590
rect 36428 20526 36430 20578
rect 36482 20526 36484 20578
rect 36428 20244 36484 20526
rect 36428 20178 36484 20188
rect 36876 20020 36932 22092
rect 36988 21700 37044 21710
rect 36988 21586 37044 21644
rect 36988 21534 36990 21586
rect 37042 21534 37044 21586
rect 36988 21522 37044 21534
rect 37212 21700 37268 21710
rect 37212 21588 37268 21644
rect 37212 21586 37380 21588
rect 37212 21534 37214 21586
rect 37266 21534 37380 21586
rect 37212 21532 37380 21534
rect 37212 21522 37268 21532
rect 37212 20802 37268 20814
rect 37212 20750 37214 20802
rect 37266 20750 37268 20802
rect 37212 20244 37268 20750
rect 37212 20178 37268 20188
rect 37100 20020 37156 20030
rect 36932 20018 37156 20020
rect 36932 19966 37102 20018
rect 37154 19966 37156 20018
rect 36932 19964 37156 19966
rect 36876 19926 36932 19964
rect 37100 19954 37156 19964
rect 37324 19906 37380 21532
rect 37324 19854 37326 19906
rect 37378 19854 37380 19906
rect 37324 19842 37380 19854
rect 37436 21364 37492 23214
rect 37660 23156 37716 23772
rect 37996 23762 38052 23772
rect 37548 23100 37716 23156
rect 38332 23380 38388 27022
rect 39564 27076 39620 27086
rect 40012 27076 40068 27086
rect 39564 27074 40068 27076
rect 39564 27022 39566 27074
rect 39618 27022 40014 27074
rect 40066 27022 40068 27074
rect 39564 27020 40068 27022
rect 39564 27010 39620 27020
rect 39564 26852 39620 26862
rect 39564 26514 39620 26796
rect 39788 26850 39844 26862
rect 39788 26798 39790 26850
rect 39842 26798 39844 26850
rect 39788 26628 39844 26798
rect 39788 26562 39844 26572
rect 39564 26462 39566 26514
rect 39618 26462 39620 26514
rect 39564 26450 39620 26462
rect 39788 26402 39844 26414
rect 39788 26350 39790 26402
rect 39842 26350 39844 26402
rect 39788 25284 39844 26350
rect 40012 26292 40068 27020
rect 40124 26852 40180 26862
rect 40124 26402 40180 26796
rect 40124 26350 40126 26402
rect 40178 26350 40180 26402
rect 40124 26338 40180 26350
rect 40012 26226 40068 26236
rect 39788 25218 39844 25228
rect 40124 24612 40180 24622
rect 40124 24518 40180 24556
rect 40124 24052 40180 24062
rect 40124 23958 40180 23996
rect 37548 21698 37604 23100
rect 37660 22932 37716 22942
rect 37660 22930 37828 22932
rect 37660 22878 37662 22930
rect 37714 22878 37828 22930
rect 37660 22876 37828 22878
rect 37660 22866 37716 22876
rect 37772 22148 37828 22876
rect 37884 22428 38276 22484
rect 37884 22370 37940 22428
rect 37884 22318 37886 22370
rect 37938 22318 37940 22370
rect 37884 22306 37940 22318
rect 38220 22370 38276 22428
rect 38220 22318 38222 22370
rect 38274 22318 38276 22370
rect 38220 22306 38276 22318
rect 37996 22258 38052 22270
rect 37996 22206 37998 22258
rect 38050 22206 38052 22258
rect 37996 22148 38052 22206
rect 37772 22092 38052 22148
rect 38332 22036 38388 23324
rect 38556 22258 38612 22270
rect 38556 22206 38558 22258
rect 38610 22206 38612 22258
rect 38444 22148 38500 22158
rect 38444 22054 38500 22092
rect 37884 21980 38388 22036
rect 37884 21810 37940 21980
rect 37884 21758 37886 21810
rect 37938 21758 37940 21810
rect 37884 21746 37940 21758
rect 37548 21646 37550 21698
rect 37602 21646 37604 21698
rect 37548 21634 37604 21646
rect 38556 21700 38612 22206
rect 38556 21634 38612 21644
rect 38108 21588 38164 21598
rect 38108 21494 38164 21532
rect 39116 21586 39172 21598
rect 39116 21534 39118 21586
rect 39170 21534 39172 21586
rect 36092 18398 36094 18450
rect 36146 18398 36148 18450
rect 35532 18338 35700 18340
rect 35532 18286 35534 18338
rect 35586 18286 35700 18338
rect 35532 18284 35700 18286
rect 35532 18274 35588 18284
rect 35308 18162 35364 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17780 35588 17790
rect 35084 17778 35588 17780
rect 35084 17726 35534 17778
rect 35586 17726 35588 17778
rect 35084 17724 35588 17726
rect 34636 16830 34638 16882
rect 34690 16830 34692 16882
rect 34636 16818 34692 16830
rect 34748 16884 34804 16894
rect 34412 16772 34468 16782
rect 34300 16770 34468 16772
rect 34300 16718 34414 16770
rect 34466 16718 34468 16770
rect 34300 16716 34468 16718
rect 34188 16706 34244 16716
rect 34412 16706 34468 16716
rect 33852 16324 33908 16334
rect 34636 16324 34692 16334
rect 33852 16322 34692 16324
rect 33852 16270 33854 16322
rect 33906 16270 34638 16322
rect 34690 16270 34692 16322
rect 33852 16268 34692 16270
rect 33852 16258 33908 16268
rect 34636 16258 34692 16268
rect 33740 15934 33742 15986
rect 33794 15934 33796 15986
rect 33740 15922 33796 15934
rect 34300 16098 34356 16110
rect 34300 16046 34302 16098
rect 34354 16046 34356 16098
rect 34300 15652 34356 16046
rect 34524 16100 34580 16110
rect 34748 16100 34804 16828
rect 34972 16882 35028 17052
rect 34972 16830 34974 16882
rect 35026 16830 35028 16882
rect 34972 16818 35028 16830
rect 35084 17444 35140 17454
rect 35084 16324 35140 17388
rect 35532 16884 35588 17724
rect 35644 17666 35700 18284
rect 36092 17892 36148 18398
rect 36540 19236 36596 19246
rect 36540 18450 36596 19180
rect 37436 19236 37492 21308
rect 37996 20690 38052 20702
rect 37996 20638 37998 20690
rect 38050 20638 38052 20690
rect 37884 19794 37940 19806
rect 37884 19742 37886 19794
rect 37938 19742 37940 19794
rect 37772 19460 37828 19470
rect 37884 19460 37940 19742
rect 37772 19458 37940 19460
rect 37772 19406 37774 19458
rect 37826 19406 37940 19458
rect 37772 19404 37940 19406
rect 37772 19394 37828 19404
rect 37996 19346 38052 20638
rect 38892 20132 38948 20142
rect 38892 20038 38948 20076
rect 39116 19796 39172 21534
rect 40124 21588 40180 21598
rect 40012 21474 40068 21486
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 20916 40068 21422
rect 40012 20850 40068 20860
rect 40124 20914 40180 21532
rect 40124 20862 40126 20914
rect 40178 20862 40180 20914
rect 40124 20850 40180 20862
rect 39676 20132 39732 20142
rect 39676 20038 39732 20076
rect 39116 19730 39172 19740
rect 37996 19294 37998 19346
rect 38050 19294 38052 19346
rect 37996 19282 38052 19294
rect 40012 19572 40068 19582
rect 40012 19346 40068 19516
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 40012 19282 40068 19294
rect 38892 19236 38948 19246
rect 37436 19142 37492 19180
rect 38556 19234 38948 19236
rect 38556 19182 38894 19234
rect 38946 19182 38948 19234
rect 38556 19180 38948 19182
rect 37100 19012 37156 19022
rect 36988 19010 37156 19012
rect 36988 18958 37102 19010
rect 37154 18958 37156 19010
rect 36988 18956 37156 18958
rect 36652 18564 36708 18574
rect 36652 18470 36708 18508
rect 36540 18398 36542 18450
rect 36594 18398 36596 18450
rect 36540 18386 36596 18398
rect 36988 18452 37044 18956
rect 37100 18946 37156 18956
rect 37996 19010 38052 19022
rect 37996 18958 37998 19010
rect 38050 18958 38052 19010
rect 37324 18676 37380 18686
rect 37324 18582 37380 18620
rect 36316 18340 36372 18350
rect 36316 18246 36372 18284
rect 36092 17826 36148 17836
rect 35644 17614 35646 17666
rect 35698 17614 35700 17666
rect 35644 17602 35700 17614
rect 36316 17556 36372 17566
rect 36316 17554 36596 17556
rect 36316 17502 36318 17554
rect 36370 17502 36596 17554
rect 36316 17500 36596 17502
rect 36316 17490 36372 17500
rect 35532 16790 35588 16828
rect 35980 17108 36036 17118
rect 35196 16772 35252 16782
rect 35196 16678 35252 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35084 16258 35140 16268
rect 34524 16098 34804 16100
rect 34524 16046 34526 16098
rect 34578 16046 34804 16098
rect 34524 16044 34804 16046
rect 34524 16034 34580 16044
rect 34300 15586 34356 15596
rect 34636 15874 34692 15886
rect 34636 15822 34638 15874
rect 34690 15822 34692 15874
rect 33404 15486 33406 15538
rect 33458 15486 33460 15538
rect 33404 15148 33460 15486
rect 33404 15092 33796 15148
rect 33404 14756 33460 14766
rect 33404 13636 33460 14700
rect 33516 14084 33572 14094
rect 33572 14028 33684 14084
rect 33516 14018 33572 14028
rect 33516 13636 33572 13646
rect 33404 13634 33572 13636
rect 33404 13582 33518 13634
rect 33570 13582 33572 13634
rect 33404 13580 33572 13582
rect 33516 13570 33572 13580
rect 33292 13122 33348 13132
rect 33180 12350 33182 12402
rect 33234 12350 33236 12402
rect 33180 12338 33236 12350
rect 33516 13074 33572 13086
rect 33516 13022 33518 13074
rect 33570 13022 33572 13074
rect 33516 12180 33572 13022
rect 33516 12114 33572 12124
rect 33628 12178 33684 14028
rect 33628 12126 33630 12178
rect 33682 12126 33684 12178
rect 33628 12114 33684 12126
rect 33740 12178 33796 15092
rect 34636 13860 34692 15822
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34636 13794 34692 13804
rect 35644 13860 35700 13870
rect 35644 13766 35700 13804
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 33740 12126 33742 12178
rect 33794 12126 33796 12178
rect 33740 12114 33796 12126
rect 33964 13188 34020 13198
rect 33964 12178 34020 13132
rect 34076 12852 34132 12862
rect 34076 12290 34132 12796
rect 35644 12852 35700 12862
rect 35644 12758 35700 12796
rect 34076 12238 34078 12290
rect 34130 12238 34132 12290
rect 34076 12226 34132 12238
rect 33964 12126 33966 12178
rect 34018 12126 34020 12178
rect 33852 11508 33908 11518
rect 33964 11508 34020 12126
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 33852 11506 34020 11508
rect 33852 11454 33854 11506
rect 33906 11454 34020 11506
rect 33852 11452 34020 11454
rect 33852 11442 33908 11452
rect 32956 11396 33012 11406
rect 32956 11302 33012 11340
rect 33516 11396 33572 11406
rect 32732 10322 32788 10332
rect 32844 11284 32900 11294
rect 32844 9940 32900 11228
rect 33292 11284 33348 11294
rect 33292 11190 33348 11228
rect 33516 10498 33572 11340
rect 33516 10446 33518 10498
rect 33570 10446 33572 10498
rect 33516 10434 33572 10446
rect 34076 10500 34132 10510
rect 32844 9846 32900 9884
rect 33852 9940 33908 9950
rect 32620 9828 32676 9838
rect 32284 9826 32676 9828
rect 32284 9774 32622 9826
rect 32674 9774 32676 9826
rect 32284 9772 32676 9774
rect 32284 9716 32340 9772
rect 32620 9762 32676 9772
rect 33852 9826 33908 9884
rect 34076 9938 34132 10444
rect 35644 10500 35700 10510
rect 35644 10406 35700 10444
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34076 9886 34078 9938
rect 34130 9886 34132 9938
rect 34076 9874 34132 9886
rect 34860 9940 34916 9950
rect 34860 9938 35252 9940
rect 34860 9886 34862 9938
rect 34914 9886 35252 9938
rect 34860 9884 35252 9886
rect 34860 9874 34916 9884
rect 33852 9774 33854 9826
rect 33906 9774 33908 9826
rect 33852 9762 33908 9774
rect 34188 9828 34244 9838
rect 34188 9734 34244 9772
rect 34748 9828 34804 9838
rect 31948 9604 32004 9614
rect 31948 9510 32004 9548
rect 31724 9102 31726 9154
rect 31778 9102 31780 9154
rect 31724 9090 31780 9102
rect 29596 8878 29598 8930
rect 29650 8878 29652 8930
rect 29596 8484 29652 8878
rect 29596 8418 29652 8428
rect 32284 8482 32340 9660
rect 33292 9716 33348 9726
rect 33292 9622 33348 9660
rect 34524 9716 34580 9726
rect 34524 9622 34580 9660
rect 34748 9714 34804 9772
rect 34748 9662 34750 9714
rect 34802 9662 34804 9714
rect 34748 9650 34804 9662
rect 32284 8430 32286 8482
rect 32338 8430 32340 8482
rect 32284 8418 32340 8430
rect 32396 9604 32452 9614
rect 32396 8370 32452 9548
rect 33068 9604 33124 9614
rect 32396 8318 32398 8370
rect 32450 8318 32452 8370
rect 32396 8306 32452 8318
rect 32508 9044 32564 9054
rect 29372 6850 29428 6860
rect 32508 8036 32564 8988
rect 33068 8930 33124 9548
rect 35196 9154 35252 9884
rect 35980 9828 36036 17052
rect 36540 16994 36596 17500
rect 36764 17108 36820 17118
rect 36988 17108 37044 18396
rect 37772 18564 37828 18574
rect 37436 18340 37492 18350
rect 37100 17668 37156 17678
rect 37100 17666 37268 17668
rect 37100 17614 37102 17666
rect 37154 17614 37268 17666
rect 37100 17612 37268 17614
rect 37100 17602 37156 17612
rect 36820 17052 37044 17108
rect 36764 17014 36820 17052
rect 36540 16942 36542 16994
rect 36594 16942 36596 16994
rect 36540 16930 36596 16942
rect 36652 16996 36708 17006
rect 36652 16902 36708 16940
rect 36204 16884 36260 16894
rect 36204 16770 36260 16828
rect 37212 16884 37268 17612
rect 37212 16790 37268 16828
rect 36204 16718 36206 16770
rect 36258 16718 36260 16770
rect 36204 15876 36260 16718
rect 37436 16212 37492 18284
rect 37772 17778 37828 18508
rect 37996 18452 38052 18958
rect 37996 18386 38052 18396
rect 38108 18228 38164 18238
rect 38108 18134 38164 18172
rect 37772 17726 37774 17778
rect 37826 17726 37828 17778
rect 37772 17714 37828 17726
rect 38556 17780 38612 19180
rect 38892 19170 38948 19180
rect 39676 18900 39732 18910
rect 38892 18452 38948 18462
rect 38892 18358 38948 18396
rect 39676 18450 39732 18844
rect 39676 18398 39678 18450
rect 39730 18398 39732 18450
rect 39676 18386 39732 18398
rect 38556 17714 38612 17724
rect 39676 17556 39732 17566
rect 37996 16996 38052 17006
rect 37996 16902 38052 16940
rect 38892 16324 38948 16334
rect 37436 16146 37492 16156
rect 38332 16212 38388 16222
rect 38332 16118 38388 16156
rect 37324 16100 37380 16110
rect 37324 16006 37380 16044
rect 38892 16098 38948 16268
rect 39676 16322 39732 17500
rect 40012 17442 40068 17454
rect 40012 17390 40014 17442
rect 40066 17390 40068 17442
rect 40012 17332 40068 17390
rect 40012 17266 40068 17276
rect 39676 16270 39678 16322
rect 39730 16270 39732 16322
rect 39676 16258 39732 16270
rect 39788 16884 39844 16894
rect 38892 16046 38894 16098
rect 38946 16046 38948 16098
rect 38892 16034 38948 16046
rect 36428 15876 36484 15886
rect 36204 15874 36484 15876
rect 36204 15822 36430 15874
rect 36482 15822 36484 15874
rect 36204 15820 36484 15822
rect 36204 14418 36260 14430
rect 36204 14366 36206 14418
rect 36258 14366 36260 14418
rect 36204 13748 36260 14366
rect 36428 13748 36484 15820
rect 37324 15876 37380 15886
rect 37324 15538 37380 15820
rect 37324 15486 37326 15538
rect 37378 15486 37380 15538
rect 37324 15474 37380 15486
rect 38892 15540 38948 15550
rect 38892 15446 38948 15484
rect 39564 15540 39620 15550
rect 38108 15202 38164 15214
rect 38108 15150 38110 15202
rect 38162 15150 38164 15202
rect 38108 14868 38164 15150
rect 38108 14802 38164 14812
rect 38892 15092 38948 15102
rect 38892 14530 38948 15036
rect 39564 14642 39620 15484
rect 39676 15540 39732 15550
rect 39788 15540 39844 16828
rect 40124 16770 40180 16782
rect 40124 16718 40126 16770
rect 40178 16718 40180 16770
rect 40124 16548 40180 16718
rect 40124 16482 40180 16492
rect 39676 15538 39844 15540
rect 39676 15486 39678 15538
rect 39730 15486 39844 15538
rect 39676 15484 39844 15486
rect 39676 15474 39732 15484
rect 39564 14590 39566 14642
rect 39618 14590 39620 14642
rect 39564 14578 39620 14590
rect 38892 14478 38894 14530
rect 38946 14478 38948 14530
rect 38892 14466 38948 14478
rect 36204 13746 36484 13748
rect 36204 13694 36430 13746
rect 36482 13694 36484 13746
rect 36204 13692 36484 13694
rect 35980 9762 36036 9772
rect 36428 13636 36484 13692
rect 36876 13636 36932 13646
rect 36428 13634 36932 13636
rect 36428 13582 36878 13634
rect 36930 13582 36932 13634
rect 36428 13580 36932 13582
rect 36428 12962 36484 13580
rect 36876 13570 36932 13580
rect 36428 12910 36430 12962
rect 36482 12910 36484 12962
rect 36428 12740 36484 12910
rect 38892 12964 38948 12974
rect 38892 12870 38948 12908
rect 40012 12852 40068 12862
rect 40012 12758 40068 12796
rect 36428 10612 36484 12684
rect 37100 12740 37156 12750
rect 37100 12646 37156 12684
rect 40124 12290 40180 12302
rect 40124 12238 40126 12290
rect 40178 12238 40180 12290
rect 40124 12180 40180 12238
rect 40124 12114 40180 12124
rect 36876 10612 36932 10622
rect 36428 10610 36932 10612
rect 36428 10558 36430 10610
rect 36482 10558 36878 10610
rect 36930 10558 36932 10610
rect 36428 10556 36932 10558
rect 35196 9102 35198 9154
rect 35250 9102 35252 9154
rect 35196 9090 35252 9102
rect 35868 9044 35924 9054
rect 35868 8950 35924 8988
rect 36428 9044 36484 10556
rect 36876 10546 36932 10556
rect 36428 8950 36484 8988
rect 33068 8878 33070 8930
rect 33122 8878 33124 8930
rect 33068 8866 33124 8878
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 38892 8260 38948 8270
rect 38668 8258 38948 8260
rect 38668 8206 38894 8258
rect 38946 8206 38948 8258
rect 38668 8204 38948 8206
rect 32844 8036 32900 8046
rect 32508 8034 32900 8036
rect 32508 7982 32846 8034
rect 32898 7982 32900 8034
rect 32508 7980 32900 7982
rect 28812 5908 28868 5918
rect 28812 5814 28868 5852
rect 32508 5908 32564 7980
rect 32844 7970 32900 7980
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 32508 5842 32564 5852
rect 38444 6020 38500 6030
rect 28364 5742 28366 5794
rect 28418 5742 28420 5794
rect 28364 5730 28420 5742
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 26124 5348 26180 5358
rect 26124 5254 26180 5292
rect 25788 5142 25844 5180
rect 26348 5236 26404 5246
rect 26404 5180 26516 5236
rect 26348 5170 26404 5180
rect 26236 5124 26292 5134
rect 26236 5030 26292 5068
rect 26460 5122 26516 5180
rect 26460 5070 26462 5122
rect 26514 5070 26516 5122
rect 26460 5058 26516 5070
rect 38444 5122 38500 5964
rect 38444 5070 38446 5122
rect 38498 5070 38500 5122
rect 38444 5058 38500 5070
rect 38668 5010 38724 8204
rect 38892 8194 38948 8204
rect 40012 8146 40068 8158
rect 40012 8094 40014 8146
rect 40066 8094 40068 8146
rect 39676 7586 39732 7598
rect 39676 7534 39678 7586
rect 39730 7534 39732 7586
rect 39676 6804 39732 7534
rect 40012 7476 40068 8094
rect 40124 8148 40180 8158
rect 40124 7698 40180 8092
rect 40124 7646 40126 7698
rect 40178 7646 40180 7698
rect 40124 7634 40180 7646
rect 40012 7410 40068 7420
rect 39676 6738 39732 6748
rect 40124 6466 40180 6478
rect 40124 6414 40126 6466
rect 40178 6414 40180 6466
rect 40124 6132 40180 6414
rect 40124 6066 40180 6076
rect 39788 6020 39844 6030
rect 39788 5926 39844 5964
rect 39564 5908 39620 5918
rect 39564 5814 39620 5852
rect 40124 5908 40180 5918
rect 40124 5460 40180 5852
rect 40124 5394 40180 5404
rect 38668 4958 38670 5010
rect 38722 4958 38724 5010
rect 38668 4946 38724 4958
rect 40124 4898 40180 4910
rect 40124 4846 40126 4898
rect 40178 4846 40180 4898
rect 40124 4788 40180 4846
rect 40124 4722 40180 4732
rect 24332 4450 24500 4452
rect 24332 4398 24334 4450
rect 24386 4398 24500 4450
rect 24332 4396 24500 4398
rect 39676 4450 39732 4462
rect 39676 4398 39678 4450
rect 39730 4398 39732 4450
rect 24332 4386 24388 4396
rect 23996 4174 23998 4226
rect 24050 4174 24052 4226
rect 23996 4162 24052 4174
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 21196 3668 21252 3678
rect 21196 3574 21252 3612
rect 20748 3556 20804 3566
rect 19852 3390 19854 3442
rect 19906 3390 19908 3442
rect 19852 3378 19908 3390
rect 20188 3444 20244 3482
rect 20748 3462 20804 3500
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 3388
rect 33180 3332 33236 3342
rect 32956 3330 33236 3332
rect 32956 3278 33182 3330
rect 33234 3278 33236 3330
rect 32956 3276 33236 3278
rect 32956 800 33012 3276
rect 33180 3266 33236 3276
rect 39228 3330 39284 3342
rect 39228 3278 39230 3330
rect 39282 3278 39284 3330
rect 39228 2100 39284 3278
rect 39676 2772 39732 4398
rect 40124 4450 40180 4462
rect 40124 4398 40126 4450
rect 40178 4398 40180 4450
rect 40124 4116 40180 4398
rect 40124 4050 40180 4060
rect 40124 3332 40180 3342
rect 40124 3238 40180 3276
rect 39676 2706 39732 2716
rect 39228 2034 39284 2044
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 32928 0 33040 800
<< via2 >>
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 38780 43036 38836 43092
rect 40124 42364 40180 42420
rect 39228 41692 39284 41748
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 39676 41074 39732 41076
rect 39676 41022 39678 41074
rect 39678 41022 39730 41074
rect 39730 41022 39732 41074
rect 39676 41020 39732 41022
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 1708 40348 1764 40404
rect 25900 40402 25956 40404
rect 25900 40350 25902 40402
rect 25902 40350 25954 40402
rect 25954 40350 25956 40402
rect 25900 40348 25956 40350
rect 26796 40348 26852 40404
rect 26572 40290 26628 40292
rect 26572 40238 26574 40290
rect 26574 40238 26626 40290
rect 26626 40238 26628 40290
rect 26572 40236 26628 40238
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4284 39676 4340 39732
rect 1708 36988 1764 37044
rect 1708 36370 1764 36372
rect 1708 36318 1710 36370
rect 1710 36318 1762 36370
rect 1762 36318 1764 36370
rect 1708 36316 1764 36318
rect 3948 26908 4004 26964
rect 1708 25116 1764 25172
rect 2044 25340 2100 25396
rect 1708 24892 1764 24948
rect 2492 24892 2548 24948
rect 2940 25116 2996 25172
rect 1932 24220 1988 24276
rect 1708 21756 1764 21812
rect 2940 24108 2996 24164
rect 4172 25004 4228 25060
rect 4172 24556 4228 24612
rect 3276 23324 3332 23380
rect 3052 21810 3108 21812
rect 3052 21758 3054 21810
rect 3054 21758 3106 21810
rect 3106 21758 3108 21810
rect 3052 21756 3108 21758
rect 1708 20188 1764 20244
rect 2380 20524 2436 20580
rect 2492 20188 2548 20244
rect 1708 19516 1764 19572
rect 2716 20018 2772 20020
rect 2716 19966 2718 20018
rect 2718 19966 2770 20018
rect 2770 19966 2772 20018
rect 2716 19964 2772 19966
rect 2492 19516 2548 19572
rect 2828 19292 2884 19348
rect 3052 19852 3108 19908
rect 3836 23324 3892 23380
rect 24220 39506 24276 39508
rect 24220 39454 24222 39506
rect 24222 39454 24274 39506
rect 24274 39454 24276 39506
rect 24220 39452 24276 39454
rect 25340 39452 25396 39508
rect 23548 39340 23604 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 8428 37772 8484 37828
rect 8204 36988 8260 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 6972 35532 7028 35588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 5628 33458 5684 33460
rect 5628 33406 5630 33458
rect 5630 33406 5682 33458
rect 5682 33406 5684 33458
rect 5628 33404 5684 33406
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5964 30268 6020 30324
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4732 28588 4788 28644
rect 6300 28642 6356 28644
rect 6300 28590 6302 28642
rect 6302 28590 6354 28642
rect 6354 28590 6356 28642
rect 6300 28588 6356 28590
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 9660 37772 9716 37828
rect 9548 37042 9604 37044
rect 9548 36990 9550 37042
rect 9550 36990 9602 37042
rect 9602 36990 9604 37042
rect 9548 36988 9604 36990
rect 9884 36540 9940 36596
rect 9772 36204 9828 36260
rect 8204 35532 8260 35588
rect 8876 35586 8932 35588
rect 8876 35534 8878 35586
rect 8878 35534 8930 35586
rect 8930 35534 8932 35586
rect 8876 35532 8932 35534
rect 10444 35756 10500 35812
rect 10780 35308 10836 35364
rect 10220 34636 10276 34692
rect 11228 35698 11284 35700
rect 11228 35646 11230 35698
rect 11230 35646 11282 35698
rect 11282 35646 11284 35698
rect 11228 35644 11284 35646
rect 7532 33180 7588 33236
rect 7644 32508 7700 32564
rect 8764 33404 8820 33460
rect 8540 33180 8596 33236
rect 9660 34130 9716 34132
rect 9660 34078 9662 34130
rect 9662 34078 9714 34130
rect 9714 34078 9716 34130
rect 9660 34076 9716 34078
rect 9212 33964 9268 34020
rect 8764 32956 8820 33012
rect 8204 32508 8260 32564
rect 8092 32396 8148 32452
rect 8652 32450 8708 32452
rect 8652 32398 8654 32450
rect 8654 32398 8706 32450
rect 8706 32398 8708 32450
rect 8652 32396 8708 32398
rect 8316 31164 8372 31220
rect 9212 31554 9268 31556
rect 9212 31502 9214 31554
rect 9214 31502 9266 31554
rect 9266 31502 9268 31554
rect 9212 31500 9268 31502
rect 8204 30322 8260 30324
rect 8204 30270 8206 30322
rect 8206 30270 8258 30322
rect 8258 30270 8260 30322
rect 8204 30268 8260 30270
rect 8876 30156 8932 30212
rect 7532 29932 7588 29988
rect 7084 29260 7140 29316
rect 6972 27244 7028 27300
rect 5628 26908 5684 26964
rect 6188 26962 6244 26964
rect 6188 26910 6190 26962
rect 6190 26910 6242 26962
rect 6242 26910 6244 26962
rect 6188 26908 6244 26910
rect 8316 29986 8372 29988
rect 8316 29934 8318 29986
rect 8318 29934 8370 29986
rect 8370 29934 8372 29986
rect 8316 29932 8372 29934
rect 8652 29426 8708 29428
rect 8652 29374 8654 29426
rect 8654 29374 8706 29426
rect 8706 29374 8708 29426
rect 8652 29372 8708 29374
rect 9660 33404 9716 33460
rect 10668 33852 10724 33908
rect 10892 34188 10948 34244
rect 10668 33628 10724 33684
rect 10108 31948 10164 32004
rect 11004 34076 11060 34132
rect 10892 34018 10948 34020
rect 10892 33966 10894 34018
rect 10894 33966 10946 34018
rect 10946 33966 10948 34018
rect 10892 33964 10948 33966
rect 10892 32956 10948 33012
rect 11340 33852 11396 33908
rect 23212 38780 23268 38836
rect 12460 37826 12516 37828
rect 12460 37774 12462 37826
rect 12462 37774 12514 37826
rect 12514 37774 12516 37826
rect 12460 37772 12516 37774
rect 12124 36594 12180 36596
rect 12124 36542 12126 36594
rect 12126 36542 12178 36594
rect 12178 36542 12180 36594
rect 12124 36540 12180 36542
rect 13356 37772 13412 37828
rect 12684 36540 12740 36596
rect 13244 37324 13300 37380
rect 12012 36482 12068 36484
rect 12012 36430 12014 36482
rect 12014 36430 12066 36482
rect 12066 36430 12068 36482
rect 12012 36428 12068 36430
rect 12684 36370 12740 36372
rect 12684 36318 12686 36370
rect 12686 36318 12738 36370
rect 12738 36318 12740 36370
rect 12684 36316 12740 36318
rect 11676 35810 11732 35812
rect 11676 35758 11678 35810
rect 11678 35758 11730 35810
rect 11730 35758 11732 35810
rect 11676 35756 11732 35758
rect 12460 36258 12516 36260
rect 12460 36206 12462 36258
rect 12462 36206 12514 36258
rect 12514 36206 12516 36258
rect 12460 36204 12516 36206
rect 12236 35644 12292 35700
rect 11676 35308 11732 35364
rect 13692 37436 13748 37492
rect 14140 37324 14196 37380
rect 13468 36988 13524 37044
rect 13804 36594 13860 36596
rect 13804 36542 13806 36594
rect 13806 36542 13858 36594
rect 13858 36542 13860 36594
rect 13804 36540 13860 36542
rect 14028 36482 14084 36484
rect 14028 36430 14030 36482
rect 14030 36430 14082 36482
rect 14082 36430 14084 36482
rect 14028 36428 14084 36430
rect 13580 36316 13636 36372
rect 13916 36258 13972 36260
rect 13916 36206 13918 36258
rect 13918 36206 13970 36258
rect 13970 36206 13972 36258
rect 13916 36204 13972 36206
rect 14812 37154 14868 37156
rect 14812 37102 14814 37154
rect 14814 37102 14866 37154
rect 14866 37102 14868 37154
rect 14812 37100 14868 37102
rect 14812 36876 14868 36932
rect 13468 35308 13524 35364
rect 11452 33180 11508 33236
rect 11564 34636 11620 34692
rect 12012 34524 12068 34580
rect 12124 34130 12180 34132
rect 12124 34078 12126 34130
rect 12126 34078 12178 34130
rect 12178 34078 12180 34130
rect 12124 34076 12180 34078
rect 11564 33628 11620 33684
rect 11452 31612 11508 31668
rect 9884 30210 9940 30212
rect 9884 30158 9886 30210
rect 9886 30158 9938 30210
rect 9938 30158 9940 30210
rect 9884 30156 9940 30158
rect 9436 29372 9492 29428
rect 9212 28754 9268 28756
rect 9212 28702 9214 28754
rect 9214 28702 9266 28754
rect 9266 28702 9268 28754
rect 9212 28700 9268 28702
rect 10108 29932 10164 29988
rect 9772 29426 9828 29428
rect 9772 29374 9774 29426
rect 9774 29374 9826 29426
rect 9826 29374 9828 29426
rect 9772 29372 9828 29374
rect 9996 29314 10052 29316
rect 9996 29262 9998 29314
rect 9998 29262 10050 29314
rect 10050 29262 10052 29314
rect 9996 29260 10052 29262
rect 10108 28924 10164 28980
rect 10332 29148 10388 29204
rect 9884 28700 9940 28756
rect 10444 28924 10500 28980
rect 9548 27858 9604 27860
rect 9548 27806 9550 27858
rect 9550 27806 9602 27858
rect 9602 27806 9604 27858
rect 9548 27804 9604 27806
rect 9436 27356 9492 27412
rect 4620 24722 4676 24724
rect 4620 24670 4622 24722
rect 4622 24670 4674 24722
rect 4674 24670 4676 24722
rect 4620 24668 4676 24670
rect 5068 25116 5124 25172
rect 6412 25004 6468 25060
rect 5292 24834 5348 24836
rect 5292 24782 5294 24834
rect 5294 24782 5346 24834
rect 5346 24782 5348 24834
rect 5292 24780 5348 24782
rect 6412 24780 6468 24836
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 8652 25228 8708 25284
rect 6300 23884 6356 23940
rect 4732 23660 4788 23716
rect 5292 23436 5348 23492
rect 5180 23324 5236 23380
rect 4396 23154 4452 23156
rect 4396 23102 4398 23154
rect 4398 23102 4450 23154
rect 4450 23102 4452 23154
rect 4396 23100 4452 23102
rect 4284 22988 4340 23044
rect 5068 23266 5124 23268
rect 5068 23214 5070 23266
rect 5070 23214 5122 23266
rect 5122 23214 5124 23266
rect 5068 23212 5124 23214
rect 4508 22876 4564 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4956 22540 5012 22596
rect 5068 22482 5124 22484
rect 5068 22430 5070 22482
rect 5070 22430 5122 22482
rect 5122 22430 5124 22482
rect 5068 22428 5124 22430
rect 4844 22204 4900 22260
rect 3500 21810 3556 21812
rect 3500 21758 3502 21810
rect 3502 21758 3554 21810
rect 3554 21758 3556 21810
rect 3500 21756 3556 21758
rect 5068 21644 5124 21700
rect 3836 21532 3892 21588
rect 5628 23154 5684 23156
rect 5628 23102 5630 23154
rect 5630 23102 5682 23154
rect 5682 23102 5684 23154
rect 5628 23100 5684 23102
rect 5628 22764 5684 22820
rect 5516 22652 5572 22708
rect 5404 22092 5460 22148
rect 4620 21586 4676 21588
rect 4620 21534 4622 21586
rect 4622 21534 4674 21586
rect 4674 21534 4676 21586
rect 4620 21532 4676 21534
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4732 20636 4788 20692
rect 3612 20524 3668 20580
rect 3164 20188 3220 20244
rect 3276 20130 3332 20132
rect 3276 20078 3278 20130
rect 3278 20078 3330 20130
rect 3330 20078 3332 20130
rect 3276 20076 3332 20078
rect 3836 20242 3892 20244
rect 3836 20190 3838 20242
rect 3838 20190 3890 20242
rect 3890 20190 3892 20242
rect 3836 20188 3892 20190
rect 3724 20130 3780 20132
rect 3724 20078 3726 20130
rect 3726 20078 3778 20130
rect 3778 20078 3780 20130
rect 3724 20076 3780 20078
rect 4172 20578 4228 20580
rect 4172 20526 4174 20578
rect 4174 20526 4226 20578
rect 4226 20526 4228 20578
rect 4172 20524 4228 20526
rect 4060 19964 4116 20020
rect 4508 20578 4564 20580
rect 4508 20526 4510 20578
rect 4510 20526 4562 20578
rect 4562 20526 4564 20578
rect 4508 20524 4564 20526
rect 1932 18396 1988 18452
rect 3612 19010 3668 19012
rect 3612 18958 3614 19010
rect 3614 18958 3666 19010
rect 3666 18958 3668 19010
rect 3612 18956 3668 18958
rect 4956 21026 5012 21028
rect 4956 20974 4958 21026
rect 4958 20974 5010 21026
rect 5010 20974 5012 21026
rect 4956 20972 5012 20974
rect 5740 21756 5796 21812
rect 5852 21644 5908 21700
rect 6524 23714 6580 23716
rect 6524 23662 6526 23714
rect 6526 23662 6578 23714
rect 6578 23662 6580 23714
rect 6524 23660 6580 23662
rect 7532 24610 7588 24612
rect 7532 24558 7534 24610
rect 7534 24558 7586 24610
rect 7586 24558 7588 24610
rect 7532 24556 7588 24558
rect 7420 23436 7476 23492
rect 6412 22764 6468 22820
rect 6524 22652 6580 22708
rect 7196 23378 7252 23380
rect 7196 23326 7198 23378
rect 7198 23326 7250 23378
rect 7250 23326 7252 23378
rect 7196 23324 7252 23326
rect 7644 23324 7700 23380
rect 9212 25282 9268 25284
rect 9212 25230 9214 25282
rect 9214 25230 9266 25282
rect 9266 25230 9268 25282
rect 9212 25228 9268 25230
rect 7980 23938 8036 23940
rect 7980 23886 7982 23938
rect 7982 23886 8034 23938
rect 8034 23886 8036 23938
rect 7980 23884 8036 23886
rect 7420 23266 7476 23268
rect 7420 23214 7422 23266
rect 7422 23214 7474 23266
rect 7474 23214 7476 23266
rect 7420 23212 7476 23214
rect 6636 22876 6692 22932
rect 6412 22540 6468 22596
rect 6300 22428 6356 22484
rect 6636 22428 6692 22484
rect 6748 22316 6804 22372
rect 6524 22146 6580 22148
rect 6524 22094 6526 22146
rect 6526 22094 6578 22146
rect 6578 22094 6580 22146
rect 6524 22092 6580 22094
rect 6748 21868 6804 21924
rect 7084 21868 7140 21924
rect 6636 21698 6692 21700
rect 6636 21646 6638 21698
rect 6638 21646 6690 21698
rect 6690 21646 6692 21698
rect 6636 21644 6692 21646
rect 6188 20972 6244 21028
rect 6748 21420 6804 21476
rect 6076 20802 6132 20804
rect 6076 20750 6078 20802
rect 6078 20750 6130 20802
rect 6130 20750 6132 20802
rect 6076 20748 6132 20750
rect 4844 20300 4900 20356
rect 4956 19964 5012 20020
rect 4732 19852 4788 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4620 19404 4676 19460
rect 4732 19346 4788 19348
rect 4732 19294 4734 19346
rect 4734 19294 4786 19346
rect 4786 19294 4788 19346
rect 4732 19292 4788 19294
rect 3724 18450 3780 18452
rect 3724 18398 3726 18450
rect 3726 18398 3778 18450
rect 3778 18398 3780 18450
rect 3724 18396 3780 18398
rect 4172 18450 4228 18452
rect 4172 18398 4174 18450
rect 4174 18398 4226 18450
rect 4226 18398 4228 18450
rect 4172 18396 4228 18398
rect 5852 20412 5908 20468
rect 5292 20130 5348 20132
rect 5292 20078 5294 20130
rect 5294 20078 5346 20130
rect 5346 20078 5348 20130
rect 5292 20076 5348 20078
rect 5292 19852 5348 19908
rect 6636 20802 6692 20804
rect 6636 20750 6638 20802
rect 6638 20750 6690 20802
rect 6690 20750 6692 20802
rect 6636 20748 6692 20750
rect 7196 21810 7252 21812
rect 7196 21758 7198 21810
rect 7198 21758 7250 21810
rect 7250 21758 7252 21810
rect 7196 21756 7252 21758
rect 7532 21698 7588 21700
rect 7532 21646 7534 21698
rect 7534 21646 7586 21698
rect 7586 21646 7588 21698
rect 7532 21644 7588 21646
rect 7196 21420 7252 21476
rect 5404 18732 5460 18788
rect 4508 18172 4564 18228
rect 5404 18172 5460 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 3612 16658 3668 16660
rect 3612 16606 3614 16658
rect 3614 16606 3666 16658
rect 3666 16606 3668 16658
rect 3612 16604 3668 16606
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4844 16380 4900 16436
rect 4956 16492 5012 16548
rect 4620 16268 4676 16324
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5068 14642 5124 14644
rect 5068 14590 5070 14642
rect 5070 14590 5122 14642
rect 5122 14590 5124 14642
rect 5068 14588 5124 14590
rect 4844 14476 4900 14532
rect 5628 17164 5684 17220
rect 5628 16492 5684 16548
rect 6188 20018 6244 20020
rect 6188 19966 6190 20018
rect 6190 19966 6242 20018
rect 6242 19966 6244 20018
rect 6188 19964 6244 19966
rect 6076 18844 6132 18900
rect 6524 19404 6580 19460
rect 8428 22316 8484 22372
rect 8652 23884 8708 23940
rect 8876 23548 8932 23604
rect 8652 22316 8708 22372
rect 8988 20860 9044 20916
rect 8540 20636 8596 20692
rect 8204 20018 8260 20020
rect 8204 19966 8206 20018
rect 8206 19966 8258 20018
rect 8258 19966 8260 20018
rect 8204 19964 8260 19966
rect 8652 20018 8708 20020
rect 8652 19966 8654 20018
rect 8654 19966 8706 20018
rect 8706 19966 8708 20018
rect 8652 19964 8708 19966
rect 6300 18956 6356 19012
rect 6412 19068 6468 19124
rect 6636 19010 6692 19012
rect 6636 18958 6638 19010
rect 6638 18958 6690 19010
rect 6690 18958 6692 19010
rect 6636 18956 6692 18958
rect 6412 18732 6468 18788
rect 6300 18562 6356 18564
rect 6300 18510 6302 18562
rect 6302 18510 6354 18562
rect 6354 18510 6356 18562
rect 6300 18508 6356 18510
rect 7196 18450 7252 18452
rect 7196 18398 7198 18450
rect 7198 18398 7250 18450
rect 7250 18398 7252 18450
rect 7196 18396 7252 18398
rect 6188 17948 6244 18004
rect 5964 17164 6020 17220
rect 6860 17948 6916 18004
rect 7532 19122 7588 19124
rect 7532 19070 7534 19122
rect 7534 19070 7586 19122
rect 7586 19070 7588 19122
rect 7532 19068 7588 19070
rect 7420 18956 7476 19012
rect 7756 19010 7812 19012
rect 7756 18958 7758 19010
rect 7758 18958 7810 19010
rect 7810 18958 7812 19010
rect 7756 18956 7812 18958
rect 7644 18562 7700 18564
rect 7644 18510 7646 18562
rect 7646 18510 7698 18562
rect 7698 18510 7700 18562
rect 7644 18508 7700 18510
rect 7532 18172 7588 18228
rect 5852 16492 5908 16548
rect 5740 16380 5796 16436
rect 6188 16322 6244 16324
rect 6188 16270 6190 16322
rect 6190 16270 6242 16322
rect 6242 16270 6244 16322
rect 6188 16268 6244 16270
rect 5964 15484 6020 15540
rect 7532 16882 7588 16884
rect 7532 16830 7534 16882
rect 7534 16830 7586 16882
rect 7586 16830 7588 16882
rect 7532 16828 7588 16830
rect 6748 16492 6804 16548
rect 7308 16156 7364 16212
rect 6412 16098 6468 16100
rect 6412 16046 6414 16098
rect 6414 16046 6466 16098
rect 6466 16046 6468 16098
rect 6412 16044 6468 16046
rect 7084 16044 7140 16100
rect 6972 15932 7028 15988
rect 5516 15314 5572 15316
rect 5516 15262 5518 15314
rect 5518 15262 5570 15314
rect 5570 15262 5572 15314
rect 5516 15260 5572 15262
rect 5516 14588 5572 14644
rect 2492 13858 2548 13860
rect 2492 13806 2494 13858
rect 2494 13806 2546 13858
rect 2546 13806 2548 13858
rect 2492 13804 2548 13806
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4844 12908 4900 12964
rect 4844 12236 4900 12292
rect 4508 12066 4564 12068
rect 4508 12014 4510 12066
rect 4510 12014 4562 12066
rect 4562 12014 4564 12066
rect 4508 12012 4564 12014
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 6972 15148 7028 15204
rect 7084 15372 7140 15428
rect 5852 14588 5908 14644
rect 5964 14530 6020 14532
rect 5964 14478 5966 14530
rect 5966 14478 6018 14530
rect 6018 14478 6020 14530
rect 5964 14476 6020 14478
rect 5852 13020 5908 13076
rect 7196 15148 7252 15204
rect 6972 14530 7028 14532
rect 6972 14478 6974 14530
rect 6974 14478 7026 14530
rect 7026 14478 7028 14530
rect 6972 14476 7028 14478
rect 6636 14418 6692 14420
rect 6636 14366 6638 14418
rect 6638 14366 6690 14418
rect 6690 14366 6692 14418
rect 6636 14364 6692 14366
rect 6188 13020 6244 13076
rect 5516 12962 5572 12964
rect 5516 12910 5518 12962
rect 5518 12910 5570 12962
rect 5570 12910 5572 12962
rect 5516 12908 5572 12910
rect 4956 12012 5012 12068
rect 2716 10780 2772 10836
rect 4956 10780 5012 10836
rect 3052 10610 3108 10612
rect 3052 10558 3054 10610
rect 3054 10558 3106 10610
rect 3106 10558 3108 10610
rect 3052 10556 3108 10558
rect 2380 10444 2436 10500
rect 4956 10444 5012 10500
rect 5740 12178 5796 12180
rect 5740 12126 5742 12178
rect 5742 12126 5794 12178
rect 5794 12126 5796 12178
rect 5740 12124 5796 12126
rect 6636 12402 6692 12404
rect 6636 12350 6638 12402
rect 6638 12350 6690 12402
rect 6690 12350 6692 12402
rect 6636 12348 6692 12350
rect 6076 12236 6132 12292
rect 5852 11676 5908 11732
rect 6748 11900 6804 11956
rect 5964 11282 6020 11284
rect 5964 11230 5966 11282
rect 5966 11230 6018 11282
rect 6018 11230 6020 11282
rect 5964 11228 6020 11230
rect 7196 11676 7252 11732
rect 6748 11228 6804 11284
rect 6300 10834 6356 10836
rect 6300 10782 6302 10834
rect 6302 10782 6354 10834
rect 6354 10782 6356 10834
rect 6300 10780 6356 10782
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 7756 16882 7812 16884
rect 7756 16830 7758 16882
rect 7758 16830 7810 16882
rect 7810 16830 7812 16882
rect 7756 16828 7812 16830
rect 7532 16604 7588 16660
rect 7644 15986 7700 15988
rect 7644 15934 7646 15986
rect 7646 15934 7698 15986
rect 7698 15934 7700 15986
rect 7644 15932 7700 15934
rect 8428 19852 8484 19908
rect 8988 19852 9044 19908
rect 8316 19234 8372 19236
rect 8316 19182 8318 19234
rect 8318 19182 8370 19234
rect 8370 19182 8372 19234
rect 8316 19180 8372 19182
rect 8988 19234 9044 19236
rect 8988 19182 8990 19234
rect 8990 19182 9042 19234
rect 9042 19182 9044 19234
rect 8988 19180 9044 19182
rect 8428 19010 8484 19012
rect 8428 18958 8430 19010
rect 8430 18958 8482 19010
rect 8482 18958 8484 19010
rect 8428 18956 8484 18958
rect 8652 18844 8708 18900
rect 8988 18844 9044 18900
rect 8428 18508 8484 18564
rect 8204 18450 8260 18452
rect 8204 18398 8206 18450
rect 8206 18398 8258 18450
rect 8258 18398 8260 18450
rect 8204 18396 8260 18398
rect 8204 18172 8260 18228
rect 8764 16882 8820 16884
rect 8764 16830 8766 16882
rect 8766 16830 8818 16882
rect 8818 16830 8820 16882
rect 8764 16828 8820 16830
rect 8092 16156 8148 16212
rect 7756 15538 7812 15540
rect 7756 15486 7758 15538
rect 7758 15486 7810 15538
rect 7810 15486 7812 15538
rect 7756 15484 7812 15486
rect 7644 15426 7700 15428
rect 7644 15374 7646 15426
rect 7646 15374 7698 15426
rect 7698 15374 7700 15426
rect 7644 15372 7700 15374
rect 7868 15314 7924 15316
rect 7868 15262 7870 15314
rect 7870 15262 7922 15314
rect 7922 15262 7924 15314
rect 7868 15260 7924 15262
rect 7420 13186 7476 13188
rect 7420 13134 7422 13186
rect 7422 13134 7474 13186
rect 7474 13134 7476 13186
rect 7420 13132 7476 13134
rect 7644 13074 7700 13076
rect 7644 13022 7646 13074
rect 7646 13022 7698 13074
rect 7698 13022 7700 13074
rect 7644 13020 7700 13022
rect 9212 20690 9268 20692
rect 9212 20638 9214 20690
rect 9214 20638 9266 20690
rect 9266 20638 9268 20690
rect 9212 20636 9268 20638
rect 10780 29148 10836 29204
rect 11116 29372 11172 29428
rect 11676 32956 11732 33012
rect 12236 33180 12292 33236
rect 11676 31948 11732 32004
rect 13580 34636 13636 34692
rect 12684 31666 12740 31668
rect 12684 31614 12686 31666
rect 12686 31614 12738 31666
rect 12738 31614 12740 31666
rect 12684 31612 12740 31614
rect 14028 35474 14084 35476
rect 14028 35422 14030 35474
rect 14030 35422 14082 35474
rect 14082 35422 14084 35474
rect 14028 35420 14084 35422
rect 15260 37436 15316 37492
rect 15484 37266 15540 37268
rect 15484 37214 15486 37266
rect 15486 37214 15538 37266
rect 15538 37214 15540 37266
rect 15484 37212 15540 37214
rect 15820 37826 15876 37828
rect 15820 37774 15822 37826
rect 15822 37774 15874 37826
rect 15874 37774 15876 37826
rect 15820 37772 15876 37774
rect 16716 37772 16772 37828
rect 15596 36988 15652 37044
rect 17612 37772 17668 37828
rect 16156 37100 16212 37156
rect 16380 37266 16436 37268
rect 16380 37214 16382 37266
rect 16382 37214 16434 37266
rect 16434 37214 16436 37266
rect 16380 37212 16436 37214
rect 15484 36428 15540 36484
rect 16044 36482 16100 36484
rect 16044 36430 16046 36482
rect 16046 36430 16098 36482
rect 16098 36430 16100 36482
rect 16044 36428 16100 36430
rect 15148 36092 15204 36148
rect 15148 34690 15204 34692
rect 15148 34638 15150 34690
rect 15150 34638 15202 34690
rect 15202 34638 15204 34690
rect 15148 34636 15204 34638
rect 14924 34524 14980 34580
rect 15260 34412 15316 34468
rect 14924 34188 14980 34244
rect 13804 33964 13860 34020
rect 14812 33404 14868 33460
rect 15484 34076 15540 34132
rect 15596 36092 15652 36148
rect 17388 37212 17444 37268
rect 16492 36988 16548 37044
rect 17276 37042 17332 37044
rect 17276 36990 17278 37042
rect 17278 36990 17330 37042
rect 17330 36990 17332 37042
rect 17276 36988 17332 36990
rect 15708 35810 15764 35812
rect 15708 35758 15710 35810
rect 15710 35758 15762 35810
rect 15762 35758 15764 35810
rect 15708 35756 15764 35758
rect 15260 33404 15316 33460
rect 16156 35420 16212 35476
rect 15708 34748 15764 34804
rect 16044 34242 16100 34244
rect 16044 34190 16046 34242
rect 16046 34190 16098 34242
rect 16098 34190 16100 34242
rect 16044 34188 16100 34190
rect 16492 35644 16548 35700
rect 16828 35644 16884 35700
rect 16268 34748 16324 34804
rect 16380 34524 16436 34580
rect 16604 34300 16660 34356
rect 16492 34242 16548 34244
rect 16492 34190 16494 34242
rect 16494 34190 16546 34242
rect 16546 34190 16548 34242
rect 16492 34188 16548 34190
rect 16604 34130 16660 34132
rect 16604 34078 16606 34130
rect 16606 34078 16658 34130
rect 16658 34078 16660 34130
rect 16604 34076 16660 34078
rect 16380 34018 16436 34020
rect 16380 33966 16382 34018
rect 16382 33966 16434 34018
rect 16434 33966 16436 34018
rect 16380 33964 16436 33966
rect 16156 33516 16212 33572
rect 12236 29372 12292 29428
rect 11676 29148 11732 29204
rect 11116 28812 11172 28868
rect 12124 28924 12180 28980
rect 11564 28642 11620 28644
rect 11564 28590 11566 28642
rect 11566 28590 11618 28642
rect 11618 28590 11620 28642
rect 11564 28588 11620 28590
rect 12012 28530 12068 28532
rect 12012 28478 12014 28530
rect 12014 28478 12066 28530
rect 12066 28478 12068 28530
rect 12012 28476 12068 28478
rect 10556 27356 10612 27412
rect 13580 29426 13636 29428
rect 13580 29374 13582 29426
rect 13582 29374 13634 29426
rect 13634 29374 13636 29426
rect 13580 29372 13636 29374
rect 12908 29314 12964 29316
rect 12908 29262 12910 29314
rect 12910 29262 12962 29314
rect 12962 29262 12964 29314
rect 12908 29260 12964 29262
rect 13916 29260 13972 29316
rect 13804 29036 13860 29092
rect 12348 28588 12404 28644
rect 12460 28812 12516 28868
rect 12572 28700 12628 28756
rect 12796 28588 12852 28644
rect 10780 25564 10836 25620
rect 10220 25394 10276 25396
rect 10220 25342 10222 25394
rect 10222 25342 10274 25394
rect 10274 25342 10276 25394
rect 10220 25340 10276 25342
rect 9772 23548 9828 23604
rect 9884 23324 9940 23380
rect 10892 25394 10948 25396
rect 10892 25342 10894 25394
rect 10894 25342 10946 25394
rect 10946 25342 10948 25394
rect 10892 25340 10948 25342
rect 11004 25282 11060 25284
rect 11004 25230 11006 25282
rect 11006 25230 11058 25282
rect 11058 25230 11060 25282
rect 11004 25228 11060 25230
rect 11452 25618 11508 25620
rect 11452 25566 11454 25618
rect 11454 25566 11506 25618
rect 11506 25566 11508 25618
rect 11452 25564 11508 25566
rect 11116 25004 11172 25060
rect 10332 24780 10388 24836
rect 10892 24780 10948 24836
rect 9548 20748 9604 20804
rect 9436 20524 9492 20580
rect 9548 20300 9604 20356
rect 9324 19628 9380 19684
rect 10108 20802 10164 20804
rect 10108 20750 10110 20802
rect 10110 20750 10162 20802
rect 10162 20750 10164 20802
rect 10108 20748 10164 20750
rect 9660 19906 9716 19908
rect 9660 19854 9662 19906
rect 9662 19854 9714 19906
rect 9714 19854 9716 19906
rect 9660 19852 9716 19854
rect 9436 19234 9492 19236
rect 9436 19182 9438 19234
rect 9438 19182 9490 19234
rect 9490 19182 9492 19234
rect 9436 19180 9492 19182
rect 9884 19180 9940 19236
rect 9660 19122 9716 19124
rect 9660 19070 9662 19122
rect 9662 19070 9714 19122
rect 9714 19070 9716 19122
rect 9660 19068 9716 19070
rect 10108 18620 10164 18676
rect 9436 18508 9492 18564
rect 10556 20300 10612 20356
rect 10892 20076 10948 20132
rect 11116 19964 11172 20020
rect 11564 24722 11620 24724
rect 11564 24670 11566 24722
rect 11566 24670 11618 24722
rect 11618 24670 11620 24722
rect 11564 24668 11620 24670
rect 12348 24610 12404 24612
rect 12348 24558 12350 24610
rect 12350 24558 12402 24610
rect 12402 24558 12404 24610
rect 12348 24556 12404 24558
rect 11564 23884 11620 23940
rect 12348 23884 12404 23940
rect 11340 22482 11396 22484
rect 11340 22430 11342 22482
rect 11342 22430 11394 22482
rect 11394 22430 11396 22482
rect 11340 22428 11396 22430
rect 11676 21756 11732 21812
rect 12012 21644 12068 21700
rect 11340 20412 11396 20468
rect 12236 20412 12292 20468
rect 12236 20018 12292 20020
rect 12236 19966 12238 20018
rect 12238 19966 12290 20018
rect 12290 19966 12292 20018
rect 12236 19964 12292 19966
rect 12124 19852 12180 19908
rect 10332 18396 10388 18452
rect 8540 16210 8596 16212
rect 8540 16158 8542 16210
rect 8542 16158 8594 16210
rect 8594 16158 8596 16210
rect 8540 16156 8596 16158
rect 8316 15484 8372 15540
rect 8204 15372 8260 15428
rect 8428 15426 8484 15428
rect 8428 15374 8430 15426
rect 8430 15374 8482 15426
rect 8482 15374 8484 15426
rect 8428 15372 8484 15374
rect 8428 14364 8484 14420
rect 8540 14028 8596 14084
rect 9100 15484 9156 15540
rect 12236 18284 12292 18340
rect 9772 15538 9828 15540
rect 9772 15486 9774 15538
rect 9774 15486 9826 15538
rect 9826 15486 9828 15538
rect 9772 15484 9828 15486
rect 8764 15314 8820 15316
rect 8764 15262 8766 15314
rect 8766 15262 8818 15314
rect 8818 15262 8820 15314
rect 8764 15260 8820 15262
rect 9772 15260 9828 15316
rect 8652 13916 8708 13972
rect 8204 13804 8260 13860
rect 8092 13356 8148 13412
rect 9436 14700 9492 14756
rect 8540 13356 8596 13412
rect 7980 12738 8036 12740
rect 7980 12686 7982 12738
rect 7982 12686 8034 12738
rect 8034 12686 8036 12738
rect 7980 12684 8036 12686
rect 7756 12124 7812 12180
rect 7532 11340 7588 11396
rect 8092 12066 8148 12068
rect 8092 12014 8094 12066
rect 8094 12014 8146 12066
rect 8146 12014 8148 12066
rect 8092 12012 8148 12014
rect 8764 12348 8820 12404
rect 8428 11394 8484 11396
rect 8428 11342 8430 11394
rect 8430 11342 8482 11394
rect 8482 11342 8484 11394
rect 8428 11340 8484 11342
rect 8316 10834 8372 10836
rect 8316 10782 8318 10834
rect 8318 10782 8370 10834
rect 8370 10782 8372 10834
rect 8316 10780 8372 10782
rect 8204 10444 8260 10500
rect 8764 11394 8820 11396
rect 8764 11342 8766 11394
rect 8766 11342 8818 11394
rect 8818 11342 8820 11394
rect 8764 11340 8820 11342
rect 8764 11170 8820 11172
rect 8764 11118 8766 11170
rect 8766 11118 8818 11170
rect 8818 11118 8820 11170
rect 8764 11116 8820 11118
rect 8988 12738 9044 12740
rect 8988 12686 8990 12738
rect 8990 12686 9042 12738
rect 9042 12686 9044 12738
rect 8988 12684 9044 12686
rect 9212 13916 9268 13972
rect 9324 13692 9380 13748
rect 11564 16380 11620 16436
rect 13468 28530 13524 28532
rect 13468 28478 13470 28530
rect 13470 28478 13522 28530
rect 13522 28478 13524 28530
rect 13468 28476 13524 28478
rect 12908 28364 12964 28420
rect 13580 28418 13636 28420
rect 13580 28366 13582 28418
rect 13582 28366 13634 28418
rect 13634 28366 13636 28418
rect 13580 28364 13636 28366
rect 12572 20018 12628 20020
rect 12572 19966 12574 20018
rect 12574 19966 12626 20018
rect 12626 19966 12628 20018
rect 12572 19964 12628 19966
rect 15148 31836 15204 31892
rect 16044 33346 16100 33348
rect 16044 33294 16046 33346
rect 16046 33294 16098 33346
rect 16098 33294 16100 33346
rect 16044 33292 16100 33294
rect 15820 32508 15876 32564
rect 15820 31890 15876 31892
rect 15820 31838 15822 31890
rect 15822 31838 15874 31890
rect 15874 31838 15876 31890
rect 15820 31836 15876 31838
rect 15932 32956 15988 33012
rect 14140 28028 14196 28084
rect 14252 26908 14308 26964
rect 16380 30828 16436 30884
rect 16156 29596 16212 29652
rect 15708 29372 15764 29428
rect 16156 29148 16212 29204
rect 16156 28588 16212 28644
rect 15932 27858 15988 27860
rect 15932 27806 15934 27858
rect 15934 27806 15986 27858
rect 15986 27806 15988 27858
rect 15932 27804 15988 27806
rect 16940 31836 16996 31892
rect 17500 35308 17556 35364
rect 21420 37938 21476 37940
rect 21420 37886 21422 37938
rect 21422 37886 21474 37938
rect 21474 37886 21476 37938
rect 21420 37884 21476 37886
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 17836 37100 17892 37156
rect 17836 36482 17892 36484
rect 17836 36430 17838 36482
rect 17838 36430 17890 36482
rect 17890 36430 17892 36482
rect 17836 36428 17892 36430
rect 19852 36988 19908 37044
rect 18060 35308 18116 35364
rect 17612 34524 17668 34580
rect 17052 33180 17108 33236
rect 16604 31778 16660 31780
rect 16604 31726 16606 31778
rect 16606 31726 16658 31778
rect 16658 31726 16660 31778
rect 16604 31724 16660 31726
rect 16716 30156 16772 30212
rect 16716 29820 16772 29876
rect 16716 29650 16772 29652
rect 16716 29598 16718 29650
rect 16718 29598 16770 29650
rect 16770 29598 16772 29650
rect 16716 29596 16772 29598
rect 16940 29484 16996 29540
rect 17164 33292 17220 33348
rect 18956 35756 19012 35812
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19404 35644 19460 35700
rect 20972 36428 21028 36484
rect 23212 37884 23268 37940
rect 22540 36988 22596 37044
rect 21756 36482 21812 36484
rect 21756 36430 21758 36482
rect 21758 36430 21810 36482
rect 21810 36430 21812 36482
rect 21756 36428 21812 36430
rect 21868 36316 21924 36372
rect 25564 39452 25620 39508
rect 25564 38834 25620 38836
rect 25564 38782 25566 38834
rect 25566 38782 25618 38834
rect 25618 38782 25620 38834
rect 25564 38780 25620 38782
rect 29148 40402 29204 40404
rect 29148 40350 29150 40402
rect 29150 40350 29202 40402
rect 29202 40350 29204 40402
rect 29148 40348 29204 40350
rect 29596 40402 29652 40404
rect 29596 40350 29598 40402
rect 29598 40350 29650 40402
rect 29650 40350 29652 40402
rect 29596 40348 29652 40350
rect 27244 40236 27300 40292
rect 27356 39506 27412 39508
rect 27356 39454 27358 39506
rect 27358 39454 27410 39506
rect 27410 39454 27412 39506
rect 27356 39452 27412 39454
rect 26796 39394 26852 39396
rect 26796 39342 26798 39394
rect 26798 39342 26850 39394
rect 26850 39342 26852 39394
rect 26796 39340 26852 39342
rect 27916 38722 27972 38724
rect 27916 38670 27918 38722
rect 27918 38670 27970 38722
rect 27970 38670 27972 38722
rect 27916 38668 27972 38670
rect 23436 36988 23492 37044
rect 19404 34802 19460 34804
rect 19404 34750 19406 34802
rect 19406 34750 19458 34802
rect 19458 34750 19460 34802
rect 19404 34748 19460 34750
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 20188 34300 20244 34356
rect 19516 34242 19572 34244
rect 19516 34190 19518 34242
rect 19518 34190 19570 34242
rect 19570 34190 19572 34242
rect 19516 34188 19572 34190
rect 19852 34188 19908 34244
rect 18620 33570 18676 33572
rect 18620 33518 18622 33570
rect 18622 33518 18674 33570
rect 18674 33518 18676 33570
rect 18620 33516 18676 33518
rect 18396 33180 18452 33236
rect 18956 32732 19012 32788
rect 17388 32562 17444 32564
rect 17388 32510 17390 32562
rect 17390 32510 17442 32562
rect 17442 32510 17444 32562
rect 17388 32508 17444 32510
rect 17724 32284 17780 32340
rect 18396 32508 18452 32564
rect 17164 31948 17220 32004
rect 16380 27858 16436 27860
rect 16380 27806 16382 27858
rect 16382 27806 16434 27858
rect 16434 27806 16436 27858
rect 16380 27804 16436 27806
rect 14140 25564 14196 25620
rect 14028 24780 14084 24836
rect 13356 24668 13412 24724
rect 14252 23772 14308 23828
rect 13020 23154 13076 23156
rect 13020 23102 13022 23154
rect 13022 23102 13074 23154
rect 13074 23102 13076 23154
rect 13020 23100 13076 23102
rect 18172 31724 18228 31780
rect 17500 30882 17556 30884
rect 17500 30830 17502 30882
rect 17502 30830 17554 30882
rect 17554 30830 17556 30882
rect 17500 30828 17556 30830
rect 16716 27132 16772 27188
rect 17500 29538 17556 29540
rect 17500 29486 17502 29538
rect 17502 29486 17554 29538
rect 17554 29486 17556 29538
rect 17500 29484 17556 29486
rect 17388 29426 17444 29428
rect 17388 29374 17390 29426
rect 17390 29374 17442 29426
rect 17442 29374 17444 29426
rect 17388 29372 17444 29374
rect 17500 29202 17556 29204
rect 17500 29150 17502 29202
rect 17502 29150 17554 29202
rect 17554 29150 17556 29202
rect 17500 29148 17556 29150
rect 17500 28812 17556 28868
rect 17948 30210 18004 30212
rect 17948 30158 17950 30210
rect 17950 30158 18002 30210
rect 18002 30158 18004 30210
rect 17948 30156 18004 30158
rect 18284 30716 18340 30772
rect 19740 34076 19796 34132
rect 19292 33516 19348 33572
rect 19516 33234 19572 33236
rect 19516 33182 19518 33234
rect 19518 33182 19570 33234
rect 19570 33182 19572 33234
rect 20300 34130 20356 34132
rect 20300 34078 20302 34130
rect 20302 34078 20354 34130
rect 20354 34078 20356 34130
rect 20300 34076 20356 34078
rect 19516 33180 19572 33182
rect 18844 32562 18900 32564
rect 18844 32510 18846 32562
rect 18846 32510 18898 32562
rect 18898 32510 18900 32562
rect 18844 32508 18900 32510
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19740 32732 19796 32788
rect 19404 32562 19460 32564
rect 19404 32510 19406 32562
rect 19406 32510 19458 32562
rect 19458 32510 19460 32562
rect 19404 32508 19460 32510
rect 19068 32284 19124 32340
rect 18508 31778 18564 31780
rect 18508 31726 18510 31778
rect 18510 31726 18562 31778
rect 18562 31726 18564 31778
rect 18508 31724 18564 31726
rect 19852 31836 19908 31892
rect 20076 31724 20132 31780
rect 20412 35644 20468 35700
rect 20524 34188 20580 34244
rect 23324 36316 23380 36372
rect 21532 33964 21588 34020
rect 20636 32732 20692 32788
rect 20636 32508 20692 32564
rect 20300 32284 20356 32340
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19068 30770 19124 30772
rect 19068 30718 19070 30770
rect 19070 30718 19122 30770
rect 19122 30718 19124 30770
rect 19068 30716 19124 30718
rect 18732 30156 18788 30212
rect 18508 29986 18564 29988
rect 18508 29934 18510 29986
rect 18510 29934 18562 29986
rect 18562 29934 18564 29986
rect 18508 29932 18564 29934
rect 18396 29596 18452 29652
rect 18060 29036 18116 29092
rect 18172 28642 18228 28644
rect 18172 28590 18174 28642
rect 18174 28590 18226 28642
rect 18226 28590 18228 28642
rect 18172 28588 18228 28590
rect 19180 29820 19236 29876
rect 19404 29932 19460 29988
rect 18844 28812 18900 28868
rect 18732 27692 18788 27748
rect 18508 27132 18564 27188
rect 16380 23714 16436 23716
rect 16380 23662 16382 23714
rect 16382 23662 16434 23714
rect 16434 23662 16436 23714
rect 16380 23660 16436 23662
rect 15484 23266 15540 23268
rect 15484 23214 15486 23266
rect 15486 23214 15538 23266
rect 15538 23214 15540 23266
rect 15484 23212 15540 23214
rect 16380 23266 16436 23268
rect 16380 23214 16382 23266
rect 16382 23214 16434 23266
rect 16434 23214 16436 23266
rect 16380 23212 16436 23214
rect 16268 23154 16324 23156
rect 16268 23102 16270 23154
rect 16270 23102 16322 23154
rect 16322 23102 16324 23154
rect 16268 23100 16324 23102
rect 15708 22540 15764 22596
rect 14476 21868 14532 21924
rect 13916 21698 13972 21700
rect 13916 21646 13918 21698
rect 13918 21646 13970 21698
rect 13970 21646 13972 21698
rect 13916 21644 13972 21646
rect 15372 21698 15428 21700
rect 15372 21646 15374 21698
rect 15374 21646 15426 21698
rect 15426 21646 15428 21698
rect 15372 21644 15428 21646
rect 16828 23884 16884 23940
rect 16828 23660 16884 23716
rect 16044 21868 16100 21924
rect 15260 21586 15316 21588
rect 15260 21534 15262 21586
rect 15262 21534 15314 21586
rect 15314 21534 15316 21586
rect 15260 21532 15316 21534
rect 15596 21474 15652 21476
rect 15596 21422 15598 21474
rect 15598 21422 15650 21474
rect 15650 21422 15652 21474
rect 15596 21420 15652 21422
rect 13580 21308 13636 21364
rect 16716 22540 16772 22596
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 16268 21308 16324 21364
rect 16716 21868 16772 21924
rect 17724 26850 17780 26852
rect 17724 26798 17726 26850
rect 17726 26798 17778 26850
rect 17778 26798 17780 26850
rect 17724 26796 17780 26798
rect 17612 26460 17668 26516
rect 18396 26460 18452 26516
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20412 29372 20468 29428
rect 19852 29148 19908 29204
rect 19628 29036 19684 29092
rect 19404 27746 19460 27748
rect 19404 27694 19406 27746
rect 19406 27694 19458 27746
rect 19458 27694 19460 27746
rect 19404 27692 19460 27694
rect 19292 27132 19348 27188
rect 18508 25004 18564 25060
rect 17052 23938 17108 23940
rect 17052 23886 17054 23938
rect 17054 23886 17106 23938
rect 17106 23886 17108 23938
rect 17052 23884 17108 23886
rect 17276 23938 17332 23940
rect 17276 23886 17278 23938
rect 17278 23886 17330 23938
rect 17330 23886 17332 23938
rect 17276 23884 17332 23886
rect 17612 24610 17668 24612
rect 17612 24558 17614 24610
rect 17614 24558 17666 24610
rect 17666 24558 17668 24610
rect 17612 24556 17668 24558
rect 17836 24108 17892 24164
rect 18508 23996 18564 24052
rect 18172 23884 18228 23940
rect 18060 23772 18116 23828
rect 17612 22540 17668 22596
rect 18172 23714 18228 23716
rect 18172 23662 18174 23714
rect 18174 23662 18226 23714
rect 18226 23662 18228 23714
rect 18172 23660 18228 23662
rect 17948 23154 18004 23156
rect 17948 23102 17950 23154
rect 17950 23102 18002 23154
rect 18002 23102 18004 23154
rect 17948 23100 18004 23102
rect 18508 23154 18564 23156
rect 18508 23102 18510 23154
rect 18510 23102 18562 23154
rect 18562 23102 18564 23154
rect 18508 23100 18564 23102
rect 17500 21756 17556 21812
rect 17052 21308 17108 21364
rect 16828 21084 16884 21140
rect 17388 21084 17444 21140
rect 13468 20412 13524 20468
rect 13804 20188 13860 20244
rect 13132 20130 13188 20132
rect 13132 20078 13134 20130
rect 13134 20078 13186 20130
rect 13186 20078 13188 20130
rect 13132 20076 13188 20078
rect 12796 19458 12852 19460
rect 12796 19406 12798 19458
rect 12798 19406 12850 19458
rect 12850 19406 12852 19458
rect 12796 19404 12852 19406
rect 12572 19234 12628 19236
rect 12572 19182 12574 19234
rect 12574 19182 12626 19234
rect 12626 19182 12628 19234
rect 12572 19180 12628 19182
rect 12796 18396 12852 18452
rect 13020 18396 13076 18452
rect 12908 18060 12964 18116
rect 12460 15484 12516 15540
rect 9660 13970 9716 13972
rect 9660 13918 9662 13970
rect 9662 13918 9714 13970
rect 9714 13918 9716 13970
rect 9660 13916 9716 13918
rect 9996 13858 10052 13860
rect 9996 13806 9998 13858
rect 9998 13806 10050 13858
rect 10050 13806 10052 13858
rect 9996 13804 10052 13806
rect 11900 15148 11956 15204
rect 12460 15036 12516 15092
rect 12348 14530 12404 14532
rect 12348 14478 12350 14530
rect 12350 14478 12402 14530
rect 12402 14478 12404 14530
rect 12348 14476 12404 14478
rect 11452 13746 11508 13748
rect 11452 13694 11454 13746
rect 11454 13694 11506 13746
rect 11506 13694 11508 13746
rect 11452 13692 11508 13694
rect 10332 13580 10388 13636
rect 11004 13580 11060 13636
rect 9660 13132 9716 13188
rect 9548 12796 9604 12852
rect 9884 12572 9940 12628
rect 9660 12066 9716 12068
rect 9660 12014 9662 12066
rect 9662 12014 9714 12066
rect 9714 12014 9716 12066
rect 9660 12012 9716 12014
rect 9436 11452 9492 11508
rect 9212 11340 9268 11396
rect 10444 12850 10500 12852
rect 10444 12798 10446 12850
rect 10446 12798 10498 12850
rect 10498 12798 10500 12850
rect 10444 12796 10500 12798
rect 9996 12402 10052 12404
rect 9996 12350 9998 12402
rect 9998 12350 10050 12402
rect 10050 12350 10052 12402
rect 9996 12348 10052 12350
rect 10668 11900 10724 11956
rect 10556 11506 10612 11508
rect 10556 11454 10558 11506
rect 10558 11454 10610 11506
rect 10610 11454 10612 11506
rect 10556 11452 10612 11454
rect 9100 11228 9156 11284
rect 10108 11282 10164 11284
rect 10108 11230 10110 11282
rect 10110 11230 10162 11282
rect 10162 11230 10164 11282
rect 10108 11228 10164 11230
rect 9772 11116 9828 11172
rect 9996 10668 10052 10724
rect 10108 10610 10164 10612
rect 10108 10558 10110 10610
rect 10110 10558 10162 10610
rect 10162 10558 10164 10610
rect 10108 10556 10164 10558
rect 10556 10722 10612 10724
rect 10556 10670 10558 10722
rect 10558 10670 10610 10722
rect 10610 10670 10612 10722
rect 10556 10668 10612 10670
rect 10332 10556 10388 10612
rect 8876 10498 8932 10500
rect 8876 10446 8878 10498
rect 8878 10446 8930 10498
rect 8930 10446 8932 10498
rect 8876 10444 8932 10446
rect 6300 8316 6356 8372
rect 8092 8316 8148 8372
rect 9436 8652 9492 8708
rect 10892 8316 10948 8372
rect 11340 13468 11396 13524
rect 12012 13468 12068 13524
rect 11564 12572 11620 12628
rect 11900 12738 11956 12740
rect 11900 12686 11902 12738
rect 11902 12686 11954 12738
rect 11954 12686 11956 12738
rect 11900 12684 11956 12686
rect 12460 13692 12516 13748
rect 12908 14252 12964 14308
rect 12572 12572 12628 12628
rect 12236 12460 12292 12516
rect 11788 12348 11844 12404
rect 13356 19852 13412 19908
rect 13468 19404 13524 19460
rect 13580 19628 13636 19684
rect 14252 20018 14308 20020
rect 14252 19966 14254 20018
rect 14254 19966 14306 20018
rect 14306 19966 14308 20018
rect 14252 19964 14308 19966
rect 14588 20130 14644 20132
rect 14588 20078 14590 20130
rect 14590 20078 14642 20130
rect 14642 20078 14644 20130
rect 14588 20076 14644 20078
rect 14476 19852 14532 19908
rect 14028 19234 14084 19236
rect 14028 19182 14030 19234
rect 14030 19182 14082 19234
rect 14082 19182 14084 19234
rect 14028 19180 14084 19182
rect 13692 18450 13748 18452
rect 13692 18398 13694 18450
rect 13694 18398 13746 18450
rect 13746 18398 13748 18450
rect 13692 18396 13748 18398
rect 13244 18284 13300 18340
rect 14252 18226 14308 18228
rect 14252 18174 14254 18226
rect 14254 18174 14306 18226
rect 14306 18174 14308 18226
rect 14252 18172 14308 18174
rect 15372 19234 15428 19236
rect 15372 19182 15374 19234
rect 15374 19182 15426 19234
rect 15426 19182 15428 19234
rect 15372 19180 15428 19182
rect 14476 17612 14532 17668
rect 13916 15484 13972 15540
rect 13468 14418 13524 14420
rect 13468 14366 13470 14418
rect 13470 14366 13522 14418
rect 13522 14366 13524 14418
rect 13468 14364 13524 14366
rect 14364 15090 14420 15092
rect 14364 15038 14366 15090
rect 14366 15038 14418 15090
rect 14418 15038 14420 15090
rect 14364 15036 14420 15038
rect 16380 20748 16436 20804
rect 16044 17612 16100 17668
rect 16828 17948 16884 18004
rect 15484 17388 15540 17444
rect 16716 17442 16772 17444
rect 16716 17390 16718 17442
rect 16718 17390 16770 17442
rect 16770 17390 16772 17442
rect 16716 17388 16772 17390
rect 16044 15484 16100 15540
rect 15036 14812 15092 14868
rect 14028 14530 14084 14532
rect 14028 14478 14030 14530
rect 14030 14478 14082 14530
rect 14082 14478 14084 14530
rect 14028 14476 14084 14478
rect 13692 14252 13748 14308
rect 13468 13970 13524 13972
rect 13468 13918 13470 13970
rect 13470 13918 13522 13970
rect 13522 13918 13524 13970
rect 13468 13916 13524 13918
rect 13356 13692 13412 13748
rect 14028 13746 14084 13748
rect 14028 13694 14030 13746
rect 14030 13694 14082 13746
rect 14082 13694 14084 13746
rect 14028 13692 14084 13694
rect 13804 13634 13860 13636
rect 13804 13582 13806 13634
rect 13806 13582 13858 13634
rect 13858 13582 13860 13634
rect 13804 13580 13860 13582
rect 15372 14812 15428 14868
rect 16380 15538 16436 15540
rect 16380 15486 16382 15538
rect 16382 15486 16434 15538
rect 16434 15486 16436 15538
rect 16380 15484 16436 15486
rect 16716 16716 16772 16772
rect 16828 16268 16884 16324
rect 17276 20802 17332 20804
rect 17276 20750 17278 20802
rect 17278 20750 17330 20802
rect 17330 20750 17332 20802
rect 17276 20748 17332 20750
rect 17164 20690 17220 20692
rect 17164 20638 17166 20690
rect 17166 20638 17218 20690
rect 17218 20638 17220 20690
rect 17164 20636 17220 20638
rect 17388 19292 17444 19348
rect 17388 18956 17444 19012
rect 17724 20972 17780 21028
rect 17052 18396 17108 18452
rect 17388 18284 17444 18340
rect 16604 15484 16660 15540
rect 15372 14418 15428 14420
rect 15372 14366 15374 14418
rect 15374 14366 15426 14418
rect 15426 14366 15428 14418
rect 15372 14364 15428 14366
rect 16156 14418 16212 14420
rect 16156 14366 16158 14418
rect 16158 14366 16210 14418
rect 16210 14366 16212 14418
rect 16156 14364 16212 14366
rect 15596 13916 15652 13972
rect 14924 13692 14980 13748
rect 14700 13634 14756 13636
rect 14700 13582 14702 13634
rect 14702 13582 14754 13634
rect 14754 13582 14756 13634
rect 14700 13580 14756 13582
rect 14252 13468 14308 13524
rect 13580 12684 13636 12740
rect 13132 12012 13188 12068
rect 13468 12460 13524 12516
rect 11228 11676 11284 11732
rect 11900 11452 11956 11508
rect 13580 12402 13636 12404
rect 13580 12350 13582 12402
rect 13582 12350 13634 12402
rect 13634 12350 13636 12402
rect 13580 12348 13636 12350
rect 15036 13468 15092 13524
rect 14028 12236 14084 12292
rect 14028 11900 14084 11956
rect 14140 12124 14196 12180
rect 14028 11676 14084 11732
rect 12908 11340 12964 11396
rect 12124 10610 12180 10612
rect 12124 10558 12126 10610
rect 12126 10558 12178 10610
rect 12178 10558 12180 10610
rect 12124 10556 12180 10558
rect 13580 11394 13636 11396
rect 13580 11342 13582 11394
rect 13582 11342 13634 11394
rect 13634 11342 13636 11394
rect 13580 11340 13636 11342
rect 11452 8370 11508 8372
rect 11452 8318 11454 8370
rect 11454 8318 11506 8370
rect 11506 8318 11508 8370
rect 11452 8316 11508 8318
rect 13132 8316 13188 8372
rect 13132 7474 13188 7476
rect 13132 7422 13134 7474
rect 13134 7422 13186 7474
rect 13186 7422 13188 7474
rect 13132 7420 13188 7422
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 15484 13634 15540 13636
rect 15484 13582 15486 13634
rect 15486 13582 15538 13634
rect 15538 13582 15540 13634
rect 15484 13580 15540 13582
rect 15932 13746 15988 13748
rect 15932 13694 15934 13746
rect 15934 13694 15986 13746
rect 15986 13694 15988 13746
rect 15932 13692 15988 13694
rect 15596 12460 15652 12516
rect 15260 12348 15316 12404
rect 15708 12178 15764 12180
rect 15708 12126 15710 12178
rect 15710 12126 15762 12178
rect 15762 12126 15764 12178
rect 15708 12124 15764 12126
rect 14588 12012 14644 12068
rect 15148 12012 15204 12068
rect 15708 11788 15764 11844
rect 15148 11506 15204 11508
rect 15148 11454 15150 11506
rect 15150 11454 15202 11506
rect 15202 11454 15204 11506
rect 15148 11452 15204 11454
rect 17052 16716 17108 16772
rect 16716 15372 16772 15428
rect 18396 21756 18452 21812
rect 17948 21644 18004 21700
rect 18172 21586 18228 21588
rect 18172 21534 18174 21586
rect 18174 21534 18226 21586
rect 18226 21534 18228 21586
rect 18172 21532 18228 21534
rect 17948 20972 18004 21028
rect 18060 21308 18116 21364
rect 17836 20802 17892 20804
rect 17836 20750 17838 20802
rect 17838 20750 17890 20802
rect 17890 20750 17892 20802
rect 17836 20748 17892 20750
rect 18172 20690 18228 20692
rect 18172 20638 18174 20690
rect 18174 20638 18226 20690
rect 18226 20638 18228 20690
rect 18172 20636 18228 20638
rect 18172 20242 18228 20244
rect 18172 20190 18174 20242
rect 18174 20190 18226 20242
rect 18226 20190 18228 20242
rect 18172 20188 18228 20190
rect 18284 19964 18340 20020
rect 18060 19740 18116 19796
rect 17836 18450 17892 18452
rect 17836 18398 17838 18450
rect 17838 18398 17890 18450
rect 17890 18398 17892 18450
rect 17836 18396 17892 18398
rect 17612 18284 17668 18340
rect 17836 17890 17892 17892
rect 17836 17838 17838 17890
rect 17838 17838 17890 17890
rect 17890 17838 17892 17890
rect 17836 17836 17892 17838
rect 18620 22428 18676 22484
rect 18732 22204 18788 22260
rect 19180 26514 19236 26516
rect 19180 26462 19182 26514
rect 19182 26462 19234 26514
rect 19234 26462 19236 26514
rect 19180 26460 19236 26462
rect 19068 26348 19124 26404
rect 18956 24050 19012 24052
rect 18956 23998 18958 24050
rect 18958 23998 19010 24050
rect 19010 23998 19012 24050
rect 18956 23996 19012 23998
rect 19404 26684 19460 26740
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20412 27074 20468 27076
rect 20412 27022 20414 27074
rect 20414 27022 20466 27074
rect 20466 27022 20468 27074
rect 20412 27020 20468 27022
rect 19628 26850 19684 26852
rect 19628 26798 19630 26850
rect 19630 26798 19682 26850
rect 19682 26798 19684 26850
rect 19628 26796 19684 26798
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19068 23042 19124 23044
rect 19068 22990 19070 23042
rect 19070 22990 19122 23042
rect 19122 22990 19124 23042
rect 19068 22988 19124 22990
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20188 24108 20244 24164
rect 19852 23938 19908 23940
rect 19852 23886 19854 23938
rect 19854 23886 19906 23938
rect 19906 23886 19908 23938
rect 19852 23884 19908 23886
rect 20188 23826 20244 23828
rect 20188 23774 20190 23826
rect 20190 23774 20242 23826
rect 20242 23774 20244 23826
rect 20188 23772 20244 23774
rect 20076 23714 20132 23716
rect 20076 23662 20078 23714
rect 20078 23662 20130 23714
rect 20130 23662 20132 23714
rect 20076 23660 20132 23662
rect 19628 23548 19684 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19516 22988 19572 23044
rect 19404 22428 19460 22484
rect 19292 21698 19348 21700
rect 19292 21646 19294 21698
rect 19294 21646 19346 21698
rect 19346 21646 19348 21698
rect 19292 21644 19348 21646
rect 18844 20914 18900 20916
rect 18844 20862 18846 20914
rect 18846 20862 18898 20914
rect 18898 20862 18900 20914
rect 18844 20860 18900 20862
rect 18620 20578 18676 20580
rect 18620 20526 18622 20578
rect 18622 20526 18674 20578
rect 18674 20526 18676 20578
rect 18620 20524 18676 20526
rect 19180 21532 19236 21588
rect 19068 21362 19124 21364
rect 19068 21310 19070 21362
rect 19070 21310 19122 21362
rect 19122 21310 19124 21362
rect 19068 21308 19124 21310
rect 19628 22370 19684 22372
rect 19628 22318 19630 22370
rect 19630 22318 19682 22370
rect 19682 22318 19684 22370
rect 19628 22316 19684 22318
rect 20748 31836 20804 31892
rect 21420 31724 21476 31780
rect 22428 31724 22484 31780
rect 20860 30098 20916 30100
rect 20860 30046 20862 30098
rect 20862 30046 20914 30098
rect 20914 30046 20916 30098
rect 20860 30044 20916 30046
rect 21084 29260 21140 29316
rect 20748 26962 20804 26964
rect 20748 26910 20750 26962
rect 20750 26910 20802 26962
rect 20802 26910 20804 26962
rect 20748 26908 20804 26910
rect 20636 24332 20692 24388
rect 20748 24108 20804 24164
rect 20524 22316 20580 22372
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20972 22316 21028 22372
rect 18956 20076 19012 20132
rect 19068 19852 19124 19908
rect 18956 18956 19012 19012
rect 18508 18508 18564 18564
rect 17948 16322 18004 16324
rect 17948 16270 17950 16322
rect 17950 16270 18002 16322
rect 18002 16270 18004 16322
rect 17948 16268 18004 16270
rect 17612 15820 17668 15876
rect 16716 14306 16772 14308
rect 16716 14254 16718 14306
rect 16718 14254 16770 14306
rect 16770 14254 16772 14306
rect 16716 14252 16772 14254
rect 16828 13692 16884 13748
rect 16716 12908 16772 12964
rect 16156 11676 16212 11732
rect 16604 12066 16660 12068
rect 16604 12014 16606 12066
rect 16606 12014 16658 12066
rect 16658 12014 16660 12066
rect 16604 12012 16660 12014
rect 17164 13356 17220 13412
rect 17388 14924 17444 14980
rect 18060 15874 18116 15876
rect 18060 15822 18062 15874
rect 18062 15822 18114 15874
rect 18114 15822 18116 15874
rect 18060 15820 18116 15822
rect 18172 15426 18228 15428
rect 18172 15374 18174 15426
rect 18174 15374 18226 15426
rect 18226 15374 18228 15426
rect 18172 15372 18228 15374
rect 18060 15090 18116 15092
rect 18060 15038 18062 15090
rect 18062 15038 18114 15090
rect 18114 15038 18116 15090
rect 18060 15036 18116 15038
rect 17948 14700 18004 14756
rect 17388 13804 17444 13860
rect 17500 14252 17556 14308
rect 16940 11676 16996 11732
rect 17948 14418 18004 14420
rect 17948 14366 17950 14418
rect 17950 14366 18002 14418
rect 18002 14366 18004 14418
rect 17948 14364 18004 14366
rect 17836 13804 17892 13860
rect 17612 13692 17668 13748
rect 16492 11564 16548 11620
rect 16828 11394 16884 11396
rect 16828 11342 16830 11394
rect 16830 11342 16882 11394
rect 16882 11342 16884 11394
rect 16828 11340 16884 11342
rect 14588 11228 14644 11284
rect 14364 8652 14420 8708
rect 13916 8316 13972 8372
rect 14028 8146 14084 8148
rect 14028 8094 14030 8146
rect 14030 8094 14082 8146
rect 14082 8094 14084 8146
rect 14028 8092 14084 8094
rect 16940 11282 16996 11284
rect 16940 11230 16942 11282
rect 16942 11230 16994 11282
rect 16994 11230 16996 11282
rect 16940 11228 16996 11230
rect 16044 11116 16100 11172
rect 17388 11170 17444 11172
rect 17388 11118 17390 11170
rect 17390 11118 17442 11170
rect 17442 11118 17444 11170
rect 17388 11116 17444 11118
rect 17052 10668 17108 10724
rect 18844 18674 18900 18676
rect 18844 18622 18846 18674
rect 18846 18622 18898 18674
rect 18898 18622 18900 18674
rect 18844 18620 18900 18622
rect 18620 17948 18676 18004
rect 19068 17890 19124 17892
rect 19068 17838 19070 17890
rect 19070 17838 19122 17890
rect 19122 17838 19124 17890
rect 19068 17836 19124 17838
rect 18508 16492 18564 16548
rect 18396 15372 18452 15428
rect 18508 16268 18564 16324
rect 19292 20130 19348 20132
rect 19292 20078 19294 20130
rect 19294 20078 19346 20130
rect 19346 20078 19348 20130
rect 19292 20076 19348 20078
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19740 20076 19796 20132
rect 19628 19852 19684 19908
rect 20412 20130 20468 20132
rect 20412 20078 20414 20130
rect 20414 20078 20466 20130
rect 20466 20078 20468 20130
rect 20412 20076 20468 20078
rect 19404 19010 19460 19012
rect 19404 18958 19406 19010
rect 19406 18958 19458 19010
rect 19458 18958 19460 19010
rect 19404 18956 19460 18958
rect 19404 18060 19460 18116
rect 19292 17948 19348 18004
rect 19068 16716 19124 16772
rect 19628 19068 19684 19124
rect 19964 19068 20020 19124
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20188 18844 20244 18900
rect 20300 18956 20356 19012
rect 20044 18788 20100 18790
rect 19740 18562 19796 18564
rect 19740 18510 19742 18562
rect 19742 18510 19794 18562
rect 19794 18510 19796 18562
rect 19740 18508 19796 18510
rect 20412 18508 20468 18564
rect 20636 20524 20692 20580
rect 20748 20188 20804 20244
rect 20972 20076 21028 20132
rect 20860 19964 20916 20020
rect 21532 31500 21588 31556
rect 22204 31164 22260 31220
rect 21868 30044 21924 30100
rect 21532 29986 21588 29988
rect 21532 29934 21534 29986
rect 21534 29934 21586 29986
rect 21586 29934 21588 29986
rect 21532 29932 21588 29934
rect 21420 29426 21476 29428
rect 21420 29374 21422 29426
rect 21422 29374 21474 29426
rect 21474 29374 21476 29426
rect 21420 29372 21476 29374
rect 21308 27186 21364 27188
rect 21308 27134 21310 27186
rect 21310 27134 21362 27186
rect 21362 27134 21364 27186
rect 21308 27132 21364 27134
rect 21196 24722 21252 24724
rect 21196 24670 21198 24722
rect 21198 24670 21250 24722
rect 21250 24670 21252 24722
rect 21196 24668 21252 24670
rect 22204 30268 22260 30324
rect 21532 25228 21588 25284
rect 21420 23884 21476 23940
rect 21308 23436 21364 23492
rect 21644 23660 21700 23716
rect 21308 23212 21364 23268
rect 21196 20524 21252 20580
rect 21532 21420 21588 21476
rect 22988 35586 23044 35588
rect 22988 35534 22990 35586
rect 22990 35534 23042 35586
rect 23042 35534 23044 35586
rect 22988 35532 23044 35534
rect 25116 37938 25172 37940
rect 25116 37886 25118 37938
rect 25118 37886 25170 37938
rect 25170 37886 25172 37938
rect 25116 37884 25172 37886
rect 25676 37100 25732 37156
rect 24668 36316 24724 36372
rect 23548 35532 23604 35588
rect 24780 35586 24836 35588
rect 24780 35534 24782 35586
rect 24782 35534 24834 35586
rect 24834 35534 24836 35586
rect 24780 35532 24836 35534
rect 23436 34636 23492 34692
rect 23100 33404 23156 33460
rect 22988 32620 23044 32676
rect 23212 32732 23268 32788
rect 24108 34130 24164 34132
rect 24108 34078 24110 34130
rect 24110 34078 24162 34130
rect 24162 34078 24164 34130
rect 24108 34076 24164 34078
rect 26572 37884 26628 37940
rect 26124 36876 26180 36932
rect 26460 36876 26516 36932
rect 26460 36594 26516 36596
rect 26460 36542 26462 36594
rect 26462 36542 26514 36594
rect 26514 36542 26516 36594
rect 26460 36540 26516 36542
rect 25788 35308 25844 35364
rect 27356 37938 27412 37940
rect 27356 37886 27358 37938
rect 27358 37886 27410 37938
rect 27410 37886 27412 37938
rect 27356 37884 27412 37886
rect 28252 38834 28308 38836
rect 28252 38782 28254 38834
rect 28254 38782 28306 38834
rect 28306 38782 28308 38834
rect 28252 38780 28308 38782
rect 27916 38050 27972 38052
rect 27916 37998 27918 38050
rect 27918 37998 27970 38050
rect 27970 37998 27972 38050
rect 27916 37996 27972 37998
rect 28588 37938 28644 37940
rect 28588 37886 28590 37938
rect 28590 37886 28642 37938
rect 28642 37886 28644 37938
rect 28588 37884 28644 37886
rect 28140 37826 28196 37828
rect 28140 37774 28142 37826
rect 28142 37774 28194 37826
rect 28194 37774 28196 37826
rect 28140 37772 28196 37774
rect 27916 37100 27972 37156
rect 27244 36204 27300 36260
rect 26796 35532 26852 35588
rect 26908 35532 26964 35588
rect 26684 35196 26740 35252
rect 23548 31836 23604 31892
rect 23324 31724 23380 31780
rect 22988 31164 23044 31220
rect 22988 30322 23044 30324
rect 22988 30270 22990 30322
rect 22990 30270 23042 30322
rect 23042 30270 23044 30322
rect 22988 30268 23044 30270
rect 24108 31778 24164 31780
rect 24108 31726 24110 31778
rect 24110 31726 24162 31778
rect 24162 31726 24164 31778
rect 24108 31724 24164 31726
rect 23548 31554 23604 31556
rect 23548 31502 23550 31554
rect 23550 31502 23602 31554
rect 23602 31502 23604 31554
rect 23548 31500 23604 31502
rect 23884 31500 23940 31556
rect 23772 30828 23828 30884
rect 24332 30994 24388 30996
rect 24332 30942 24334 30994
rect 24334 30942 24386 30994
rect 24386 30942 24388 30994
rect 24332 30940 24388 30942
rect 24108 30268 24164 30324
rect 22764 29932 22820 29988
rect 23324 29484 23380 29540
rect 21868 29260 21924 29316
rect 23660 28364 23716 28420
rect 22540 27244 22596 27300
rect 23324 27804 23380 27860
rect 22764 25394 22820 25396
rect 22764 25342 22766 25394
rect 22766 25342 22818 25394
rect 22818 25342 22820 25394
rect 22764 25340 22820 25342
rect 23212 25340 23268 25396
rect 22316 24834 22372 24836
rect 22316 24782 22318 24834
rect 22318 24782 22370 24834
rect 22370 24782 22372 24834
rect 22316 24780 22372 24782
rect 22092 24722 22148 24724
rect 22092 24670 22094 24722
rect 22094 24670 22146 24722
rect 22146 24670 22148 24722
rect 22092 24668 22148 24670
rect 21868 23324 21924 23380
rect 23100 23938 23156 23940
rect 23100 23886 23102 23938
rect 23102 23886 23154 23938
rect 23154 23886 23156 23938
rect 23100 23884 23156 23886
rect 22316 23660 22372 23716
rect 22764 23826 22820 23828
rect 22764 23774 22766 23826
rect 22766 23774 22818 23826
rect 22818 23774 22820 23826
rect 22764 23772 22820 23774
rect 22092 23100 22148 23156
rect 23100 23324 23156 23380
rect 23548 27020 23604 27076
rect 23436 26962 23492 26964
rect 23436 26910 23438 26962
rect 23438 26910 23490 26962
rect 23490 26910 23492 26962
rect 23436 26908 23492 26910
rect 25452 34076 25508 34132
rect 25116 33404 25172 33460
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 24668 31612 24724 31668
rect 25340 31666 25396 31668
rect 25340 31614 25342 31666
rect 25342 31614 25394 31666
rect 25394 31614 25396 31666
rect 25340 31612 25396 31614
rect 25004 31554 25060 31556
rect 25004 31502 25006 31554
rect 25006 31502 25058 31554
rect 25058 31502 25060 31554
rect 25004 31500 25060 31502
rect 24668 30492 24724 30548
rect 24556 30268 24612 30324
rect 25116 29484 25172 29540
rect 24668 28700 24724 28756
rect 24108 28252 24164 28308
rect 23772 27356 23828 27412
rect 24332 27356 24388 27412
rect 24780 28364 24836 28420
rect 24108 27020 24164 27076
rect 23884 25452 23940 25508
rect 23772 25394 23828 25396
rect 23772 25342 23774 25394
rect 23774 25342 23826 25394
rect 23826 25342 23828 25394
rect 23772 25340 23828 25342
rect 23772 23996 23828 24052
rect 24332 26572 24388 26628
rect 24780 25506 24836 25508
rect 24780 25454 24782 25506
rect 24782 25454 24834 25506
rect 24834 25454 24836 25506
rect 24780 25452 24836 25454
rect 24220 25394 24276 25396
rect 24220 25342 24222 25394
rect 24222 25342 24274 25394
rect 24274 25342 24276 25394
rect 24220 25340 24276 25342
rect 25004 24668 25060 24724
rect 22092 21868 22148 21924
rect 23100 21868 23156 21924
rect 21756 20802 21812 20804
rect 21756 20750 21758 20802
rect 21758 20750 21810 20802
rect 21810 20750 21812 20802
rect 21756 20748 21812 20750
rect 21644 20188 21700 20244
rect 20524 18396 20580 18452
rect 19628 17836 19684 17892
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 18508 14924 18564 14980
rect 18732 16156 18788 16212
rect 19516 16044 19572 16100
rect 19292 15874 19348 15876
rect 19292 15822 19294 15874
rect 19294 15822 19346 15874
rect 19346 15822 19348 15874
rect 19292 15820 19348 15822
rect 19068 15314 19124 15316
rect 19068 15262 19070 15314
rect 19070 15262 19122 15314
rect 19122 15262 19124 15314
rect 19068 15260 19124 15262
rect 18396 14812 18452 14868
rect 18956 14924 19012 14980
rect 18956 14700 19012 14756
rect 18396 14252 18452 14308
rect 19292 14364 19348 14420
rect 18284 13970 18340 13972
rect 18284 13918 18286 13970
rect 18286 13918 18338 13970
rect 18338 13918 18340 13970
rect 18284 13916 18340 13918
rect 18172 13468 18228 13524
rect 18060 13356 18116 13412
rect 17948 13244 18004 13300
rect 17836 12178 17892 12180
rect 17836 12126 17838 12178
rect 17838 12126 17890 12178
rect 17890 12126 17892 12178
rect 17836 12124 17892 12126
rect 17836 11788 17892 11844
rect 17612 11618 17668 11620
rect 17612 11566 17614 11618
rect 17614 11566 17666 11618
rect 17666 11566 17668 11618
rect 17612 11564 17668 11566
rect 17836 11394 17892 11396
rect 17836 11342 17838 11394
rect 17838 11342 17890 11394
rect 17890 11342 17892 11394
rect 17836 11340 17892 11342
rect 18956 13580 19012 13636
rect 19068 13916 19124 13972
rect 19180 13858 19236 13860
rect 19180 13806 19182 13858
rect 19182 13806 19234 13858
rect 19234 13806 19236 13858
rect 19180 13804 19236 13806
rect 20076 15932 20132 15988
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19740 15538 19796 15540
rect 19740 15486 19742 15538
rect 19742 15486 19794 15538
rect 19794 15486 19796 15538
rect 19740 15484 19796 15486
rect 19628 15314 19684 15316
rect 19628 15262 19630 15314
rect 19630 15262 19682 15314
rect 19682 15262 19684 15314
rect 19628 15260 19684 15262
rect 19740 14418 19796 14420
rect 19740 14366 19742 14418
rect 19742 14366 19794 14418
rect 19794 14366 19796 14418
rect 19740 14364 19796 14366
rect 19964 14924 20020 14980
rect 21756 20076 21812 20132
rect 21644 19404 21700 19460
rect 20972 18674 21028 18676
rect 20972 18622 20974 18674
rect 20974 18622 21026 18674
rect 21026 18622 21028 18674
rect 20972 18620 21028 18622
rect 20748 14812 20804 14868
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20300 14028 20356 14084
rect 19516 13468 19572 13524
rect 20748 14140 20804 14196
rect 20748 13970 20804 13972
rect 20748 13918 20750 13970
rect 20750 13918 20802 13970
rect 20802 13918 20804 13970
rect 20748 13916 20804 13918
rect 18956 12402 19012 12404
rect 18956 12350 18958 12402
rect 18958 12350 19010 12402
rect 19010 12350 19012 12402
rect 18956 12348 19012 12350
rect 18508 12012 18564 12068
rect 18732 11788 18788 11844
rect 18172 11676 18228 11732
rect 17948 11228 18004 11284
rect 14700 8092 14756 8148
rect 14364 7756 14420 7812
rect 15372 8428 15428 8484
rect 16380 8428 16436 8484
rect 19404 12124 19460 12180
rect 19516 12572 19572 12628
rect 19292 12012 19348 12068
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19740 12236 19796 12292
rect 21532 17724 21588 17780
rect 22316 16156 22372 16212
rect 22092 15484 22148 15540
rect 22876 16210 22932 16212
rect 22876 16158 22878 16210
rect 22878 16158 22930 16210
rect 22930 16158 22932 16210
rect 22876 16156 22932 16158
rect 23100 15596 23156 15652
rect 23772 21420 23828 21476
rect 24220 23938 24276 23940
rect 24220 23886 24222 23938
rect 24222 23886 24274 23938
rect 24274 23886 24276 23938
rect 24220 23884 24276 23886
rect 24444 23212 24500 23268
rect 25228 28700 25284 28756
rect 25788 32562 25844 32564
rect 25788 32510 25790 32562
rect 25790 32510 25842 32562
rect 25842 32510 25844 32562
rect 25788 32508 25844 32510
rect 25564 32396 25620 32452
rect 26012 32786 26068 32788
rect 26012 32734 26014 32786
rect 26014 32734 26066 32786
rect 26066 32734 26068 32786
rect 26012 32732 26068 32734
rect 26236 34076 26292 34132
rect 26012 32396 26068 32452
rect 25452 28252 25508 28308
rect 25340 27356 25396 27412
rect 25676 30940 25732 30996
rect 25788 30156 25844 30212
rect 26012 30716 26068 30772
rect 25788 28252 25844 28308
rect 25564 24780 25620 24836
rect 25788 24722 25844 24724
rect 25788 24670 25790 24722
rect 25790 24670 25842 24722
rect 25842 24670 25844 24722
rect 25788 24668 25844 24670
rect 28476 36204 28532 36260
rect 27692 35196 27748 35252
rect 26236 31724 26292 31780
rect 26572 31778 26628 31780
rect 26572 31726 26574 31778
rect 26574 31726 26626 31778
rect 26626 31726 26628 31778
rect 26572 31724 26628 31726
rect 26236 31276 26292 31332
rect 26796 31554 26852 31556
rect 26796 31502 26798 31554
rect 26798 31502 26850 31554
rect 26850 31502 26852 31554
rect 26796 31500 26852 31502
rect 27356 32786 27412 32788
rect 27356 32734 27358 32786
rect 27358 32734 27410 32786
rect 27410 32734 27412 32786
rect 27356 32732 27412 32734
rect 27020 31836 27076 31892
rect 26236 31106 26292 31108
rect 26236 31054 26238 31106
rect 26238 31054 26290 31106
rect 26290 31054 26292 31106
rect 26236 31052 26292 31054
rect 26572 30770 26628 30772
rect 26572 30718 26574 30770
rect 26574 30718 26626 30770
rect 26626 30718 26628 30770
rect 26572 30716 26628 30718
rect 26572 30492 26628 30548
rect 26460 30210 26516 30212
rect 26460 30158 26462 30210
rect 26462 30158 26514 30210
rect 26514 30158 26516 30210
rect 26460 30156 26516 30158
rect 26796 30156 26852 30212
rect 26908 30098 26964 30100
rect 26908 30046 26910 30098
rect 26910 30046 26962 30098
rect 26962 30046 26964 30098
rect 26908 30044 26964 30046
rect 27580 31836 27636 31892
rect 27132 30210 27188 30212
rect 27132 30158 27134 30210
rect 27134 30158 27186 30210
rect 27186 30158 27188 30210
rect 27132 30156 27188 30158
rect 27132 29932 27188 29988
rect 26572 29372 26628 29428
rect 27020 29538 27076 29540
rect 27020 29486 27022 29538
rect 27022 29486 27074 29538
rect 27074 29486 27076 29538
rect 27020 29484 27076 29486
rect 26908 28476 26964 28532
rect 29820 39340 29876 39396
rect 30156 38780 30212 38836
rect 29932 38668 29988 38724
rect 30156 38162 30212 38164
rect 30156 38110 30158 38162
rect 30158 38110 30210 38162
rect 30210 38110 30212 38162
rect 30156 38108 30212 38110
rect 30380 40290 30436 40292
rect 30380 40238 30382 40290
rect 30382 40238 30434 40290
rect 30434 40238 30436 40290
rect 30380 40236 30436 40238
rect 31948 40236 32004 40292
rect 30268 38556 30324 38612
rect 29148 37772 29204 37828
rect 29148 37212 29204 37268
rect 29708 37884 29764 37940
rect 29148 36540 29204 36596
rect 30268 37772 30324 37828
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 40348 40348 40404 40404
rect 40124 39676 40180 39732
rect 31276 39394 31332 39396
rect 31276 39342 31278 39394
rect 31278 39342 31330 39394
rect 31330 39342 31332 39394
rect 31276 39340 31332 39342
rect 30940 38892 30996 38948
rect 30828 37996 30884 38052
rect 31052 38108 31108 38164
rect 30492 37938 30548 37940
rect 30492 37886 30494 37938
rect 30494 37886 30546 37938
rect 30546 37886 30548 37938
rect 30492 37884 30548 37886
rect 30604 37826 30660 37828
rect 30604 37774 30606 37826
rect 30606 37774 30658 37826
rect 30658 37774 30660 37826
rect 30604 37772 30660 37774
rect 30380 37378 30436 37380
rect 30380 37326 30382 37378
rect 30382 37326 30434 37378
rect 30434 37326 30436 37378
rect 30380 37324 30436 37326
rect 30268 37266 30324 37268
rect 30268 37214 30270 37266
rect 30270 37214 30322 37266
rect 30322 37214 30324 37266
rect 30268 37212 30324 37214
rect 32060 39506 32116 39508
rect 32060 39454 32062 39506
rect 32062 39454 32114 39506
rect 32114 39454 32116 39506
rect 32060 39452 32116 39454
rect 32060 38946 32116 38948
rect 32060 38894 32062 38946
rect 32062 38894 32114 38946
rect 32114 38894 32116 38946
rect 32060 38892 32116 38894
rect 32732 38892 32788 38948
rect 31724 38668 31780 38724
rect 31612 38556 31668 38612
rect 31500 38444 31556 38500
rect 31500 37324 31556 37380
rect 31052 37212 31108 37268
rect 29708 36540 29764 36596
rect 28588 34636 28644 34692
rect 29260 34076 29316 34132
rect 28476 33458 28532 33460
rect 28476 33406 28478 33458
rect 28478 33406 28530 33458
rect 28530 33406 28532 33458
rect 28476 33404 28532 33406
rect 27916 33180 27972 33236
rect 28924 32956 28980 33012
rect 28140 32732 28196 32788
rect 27804 31836 27860 31892
rect 29036 32562 29092 32564
rect 29036 32510 29038 32562
rect 29038 32510 29090 32562
rect 29090 32510 29092 32562
rect 29036 32508 29092 32510
rect 28028 31500 28084 31556
rect 27356 27970 27412 27972
rect 27356 27918 27358 27970
rect 27358 27918 27410 27970
rect 27410 27918 27412 27970
rect 27356 27916 27412 27918
rect 27244 27804 27300 27860
rect 28364 30492 28420 30548
rect 28252 30044 28308 30100
rect 27916 28476 27972 28532
rect 27916 27804 27972 27860
rect 30380 36204 30436 36260
rect 31388 36988 31444 37044
rect 31724 37266 31780 37268
rect 31724 37214 31726 37266
rect 31726 37214 31778 37266
rect 31778 37214 31780 37266
rect 31724 37212 31780 37214
rect 31276 36258 31332 36260
rect 31276 36206 31278 36258
rect 31278 36206 31330 36258
rect 31330 36206 31332 36258
rect 31276 36204 31332 36206
rect 31500 35810 31556 35812
rect 31500 35758 31502 35810
rect 31502 35758 31554 35810
rect 31554 35758 31556 35810
rect 31500 35756 31556 35758
rect 31276 35698 31332 35700
rect 31276 35646 31278 35698
rect 31278 35646 31330 35698
rect 31330 35646 31332 35698
rect 31276 35644 31332 35646
rect 31052 35084 31108 35140
rect 31164 35420 31220 35476
rect 30492 34802 30548 34804
rect 30492 34750 30494 34802
rect 30494 34750 30546 34802
rect 30546 34750 30548 34802
rect 30492 34748 30548 34750
rect 31164 34748 31220 34804
rect 29932 34690 29988 34692
rect 29932 34638 29934 34690
rect 29934 34638 29986 34690
rect 29986 34638 29988 34690
rect 29932 34636 29988 34638
rect 29260 32562 29316 32564
rect 29260 32510 29262 32562
rect 29262 32510 29314 32562
rect 29314 32510 29316 32562
rect 29260 32508 29316 32510
rect 29708 33292 29764 33348
rect 30156 34524 30212 34580
rect 30156 34130 30212 34132
rect 30156 34078 30158 34130
rect 30158 34078 30210 34130
rect 30210 34078 30212 34130
rect 30156 34076 30212 34078
rect 30492 34354 30548 34356
rect 30492 34302 30494 34354
rect 30494 34302 30546 34354
rect 30546 34302 30548 34354
rect 30492 34300 30548 34302
rect 31052 34300 31108 34356
rect 30380 33516 30436 33572
rect 30492 34076 30548 34132
rect 30156 33404 30212 33460
rect 30380 33346 30436 33348
rect 30380 33294 30382 33346
rect 30382 33294 30434 33346
rect 30434 33294 30436 33346
rect 30380 33292 30436 33294
rect 29484 33068 29540 33124
rect 29596 31836 29652 31892
rect 30044 32284 30100 32340
rect 29484 30492 29540 30548
rect 28476 29596 28532 29652
rect 29148 29932 29204 29988
rect 29596 30044 29652 30100
rect 29260 29820 29316 29876
rect 28476 28754 28532 28756
rect 28476 28702 28478 28754
rect 28478 28702 28530 28754
rect 28530 28702 28532 28754
rect 28476 28700 28532 28702
rect 27580 26908 27636 26964
rect 27692 26290 27748 26292
rect 27692 26238 27694 26290
rect 27694 26238 27746 26290
rect 27746 26238 27748 26290
rect 27692 26236 27748 26238
rect 26236 26124 26292 26180
rect 26908 26178 26964 26180
rect 26908 26126 26910 26178
rect 26910 26126 26962 26178
rect 26962 26126 26964 26178
rect 26908 26124 26964 26126
rect 28364 26796 28420 26852
rect 28252 26124 28308 26180
rect 26684 24722 26740 24724
rect 26684 24670 26686 24722
rect 26686 24670 26738 24722
rect 26738 24670 26740 24722
rect 26684 24668 26740 24670
rect 25228 23996 25284 24052
rect 24220 21474 24276 21476
rect 24220 21422 24222 21474
rect 24222 21422 24274 21474
rect 24274 21422 24276 21474
rect 24220 21420 24276 21422
rect 23884 20748 23940 20804
rect 24668 19516 24724 19572
rect 23772 19458 23828 19460
rect 23772 19406 23774 19458
rect 23774 19406 23826 19458
rect 23826 19406 23828 19458
rect 23772 19404 23828 19406
rect 23660 19180 23716 19236
rect 24332 19234 24388 19236
rect 24332 19182 24334 19234
rect 24334 19182 24386 19234
rect 24386 19182 24388 19234
rect 24332 19180 24388 19182
rect 24780 18396 24836 18452
rect 23884 18060 23940 18116
rect 25340 21420 25396 21476
rect 25228 19906 25284 19908
rect 25228 19854 25230 19906
rect 25230 19854 25282 19906
rect 25282 19854 25284 19906
rect 25228 19852 25284 19854
rect 24892 18172 24948 18228
rect 25116 18284 25172 18340
rect 24332 18060 24388 18116
rect 24556 17778 24612 17780
rect 24556 17726 24558 17778
rect 24558 17726 24610 17778
rect 24610 17726 24612 17778
rect 24556 17724 24612 17726
rect 26348 22092 26404 22148
rect 25788 21420 25844 21476
rect 26124 21474 26180 21476
rect 26124 21422 26126 21474
rect 26126 21422 26178 21474
rect 26178 21422 26180 21474
rect 26124 21420 26180 21422
rect 27804 23436 27860 23492
rect 27468 23212 27524 23268
rect 27468 22540 27524 22596
rect 27804 22988 27860 23044
rect 26796 21756 26852 21812
rect 26908 22092 26964 22148
rect 27244 22146 27300 22148
rect 27244 22094 27246 22146
rect 27246 22094 27298 22146
rect 27298 22094 27300 22146
rect 27244 22092 27300 22094
rect 28028 22258 28084 22260
rect 28028 22206 28030 22258
rect 28030 22206 28082 22258
rect 28082 22206 28084 22258
rect 28028 22204 28084 22206
rect 27916 22092 27972 22148
rect 29036 27804 29092 27860
rect 29596 27074 29652 27076
rect 29596 27022 29598 27074
rect 29598 27022 29650 27074
rect 29650 27022 29652 27074
rect 29596 27020 29652 27022
rect 28588 26962 28644 26964
rect 28588 26910 28590 26962
rect 28590 26910 28642 26962
rect 28642 26910 28644 26962
rect 28588 26908 28644 26910
rect 29820 31554 29876 31556
rect 29820 31502 29822 31554
rect 29822 31502 29874 31554
rect 29874 31502 29876 31554
rect 29820 31500 29876 31502
rect 30156 31612 30212 31668
rect 30268 33180 30324 33236
rect 30940 34130 30996 34132
rect 30940 34078 30942 34130
rect 30942 34078 30994 34130
rect 30994 34078 30996 34130
rect 30940 34076 30996 34078
rect 31276 34690 31332 34692
rect 31276 34638 31278 34690
rect 31278 34638 31330 34690
rect 31330 34638 31332 34690
rect 31276 34636 31332 34638
rect 31276 34354 31332 34356
rect 31276 34302 31278 34354
rect 31278 34302 31330 34354
rect 31330 34302 31332 34354
rect 31276 34300 31332 34302
rect 31612 33180 31668 33236
rect 31276 33122 31332 33124
rect 31276 33070 31278 33122
rect 31278 33070 31330 33122
rect 31330 33070 31332 33122
rect 31276 33068 31332 33070
rect 31164 32956 31220 33012
rect 30828 32172 30884 32228
rect 30156 31052 30212 31108
rect 30044 30044 30100 30100
rect 30380 30098 30436 30100
rect 30380 30046 30382 30098
rect 30382 30046 30434 30098
rect 30434 30046 30436 30098
rect 30380 30044 30436 30046
rect 30268 29932 30324 29988
rect 30604 30268 30660 30324
rect 30716 30828 30772 30884
rect 31164 30492 31220 30548
rect 30828 30268 30884 30324
rect 30380 29820 30436 29876
rect 30604 29708 30660 29764
rect 30492 29596 30548 29652
rect 30268 28700 30324 28756
rect 29820 27580 29876 27636
rect 30044 27132 30100 27188
rect 28252 22428 28308 22484
rect 28588 26012 28644 26068
rect 27580 21586 27636 21588
rect 27580 21534 27582 21586
rect 27582 21534 27634 21586
rect 27634 21534 27636 21586
rect 27580 21532 27636 21534
rect 26572 21420 26628 21476
rect 25788 20748 25844 20804
rect 25900 19852 25956 19908
rect 25228 19234 25284 19236
rect 25228 19182 25230 19234
rect 25230 19182 25282 19234
rect 25282 19182 25284 19234
rect 25228 19180 25284 19182
rect 23212 17388 23268 17444
rect 21420 14812 21476 14868
rect 22764 14530 22820 14532
rect 22764 14478 22766 14530
rect 22766 14478 22818 14530
rect 22818 14478 22820 14530
rect 22764 14476 22820 14478
rect 22204 13916 22260 13972
rect 21308 13356 21364 13412
rect 21868 13356 21924 13412
rect 21196 12962 21252 12964
rect 21196 12910 21198 12962
rect 21198 12910 21250 12962
rect 21250 12910 21252 12962
rect 21196 12908 21252 12910
rect 20300 12236 20356 12292
rect 20636 12290 20692 12292
rect 20636 12238 20638 12290
rect 20638 12238 20690 12290
rect 20690 12238 20692 12290
rect 20636 12236 20692 12238
rect 20188 11452 20244 11508
rect 20076 11228 20132 11284
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19292 9996 19348 10052
rect 18172 9660 18228 9716
rect 19068 9714 19124 9716
rect 19068 9662 19070 9714
rect 19070 9662 19122 9714
rect 19122 9662 19124 9714
rect 19068 9660 19124 9662
rect 19180 9548 19236 9604
rect 18956 9154 19012 9156
rect 18956 9102 18958 9154
rect 18958 9102 19010 9154
rect 19010 9102 19012 9154
rect 18956 9100 19012 9102
rect 18844 8428 18900 8484
rect 16044 8092 16100 8148
rect 15036 7756 15092 7812
rect 14924 7644 14980 7700
rect 16044 7644 16100 7700
rect 16492 7474 16548 7476
rect 16492 7422 16494 7474
rect 16494 7422 16546 7474
rect 16546 7422 16548 7474
rect 16492 7420 16548 7422
rect 13356 6524 13412 6580
rect 1708 6466 1764 6468
rect 1708 6414 1710 6466
rect 1710 6414 1762 6466
rect 1762 6414 1764 6466
rect 1708 6412 1764 6414
rect 19068 8316 19124 8372
rect 19292 8092 19348 8148
rect 19964 10668 20020 10724
rect 19740 9996 19796 10052
rect 20412 10108 20468 10164
rect 20524 11452 20580 11508
rect 21084 11452 21140 11508
rect 21308 11282 21364 11284
rect 21308 11230 21310 11282
rect 21310 11230 21362 11282
rect 21362 11230 21364 11282
rect 21308 11228 21364 11230
rect 20748 9938 20804 9940
rect 20748 9886 20750 9938
rect 20750 9886 20802 9938
rect 20802 9886 20804 9938
rect 20748 9884 20804 9886
rect 20076 9602 20132 9604
rect 20076 9550 20078 9602
rect 20078 9550 20130 9602
rect 20130 9550 20132 9602
rect 20076 9548 20132 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20524 9772 20580 9828
rect 21420 10108 21476 10164
rect 25340 18450 25396 18452
rect 25340 18398 25342 18450
rect 25342 18398 25394 18450
rect 25394 18398 25396 18450
rect 25340 18396 25396 18398
rect 25564 18284 25620 18340
rect 25228 17724 25284 17780
rect 25564 17724 25620 17780
rect 25004 16156 25060 16212
rect 25116 16098 25172 16100
rect 25116 16046 25118 16098
rect 25118 16046 25170 16098
rect 25170 16046 25172 16098
rect 25116 16044 25172 16046
rect 25676 16044 25732 16100
rect 23436 15986 23492 15988
rect 23436 15934 23438 15986
rect 23438 15934 23490 15986
rect 23490 15934 23492 15986
rect 23436 15932 23492 15934
rect 24332 15986 24388 15988
rect 24332 15934 24334 15986
rect 24334 15934 24386 15986
rect 24386 15934 24388 15986
rect 24332 15932 24388 15934
rect 23884 15148 23940 15204
rect 23324 14476 23380 14532
rect 23772 14530 23828 14532
rect 23772 14478 23774 14530
rect 23774 14478 23826 14530
rect 23826 14478 23828 14530
rect 23772 14476 23828 14478
rect 23996 14530 24052 14532
rect 23996 14478 23998 14530
rect 23998 14478 24050 14530
rect 24050 14478 24052 14530
rect 23996 14476 24052 14478
rect 23436 14028 23492 14084
rect 24780 15932 24836 15988
rect 25340 15202 25396 15204
rect 25340 15150 25342 15202
rect 25342 15150 25394 15202
rect 25394 15150 25396 15202
rect 25340 15148 25396 15150
rect 26684 20018 26740 20020
rect 26684 19966 26686 20018
rect 26686 19966 26738 20018
rect 26738 19966 26740 20018
rect 26684 19964 26740 19966
rect 26348 19740 26404 19796
rect 26460 19906 26516 19908
rect 26460 19854 26462 19906
rect 26462 19854 26514 19906
rect 26514 19854 26516 19906
rect 26460 19852 26516 19854
rect 26236 19404 26292 19460
rect 26572 19404 26628 19460
rect 26684 18396 26740 18452
rect 26684 17442 26740 17444
rect 26684 17390 26686 17442
rect 26686 17390 26738 17442
rect 26738 17390 26740 17442
rect 26684 17388 26740 17390
rect 25116 14530 25172 14532
rect 25116 14478 25118 14530
rect 25118 14478 25170 14530
rect 25170 14478 25172 14530
rect 25116 14476 25172 14478
rect 24668 13916 24724 13972
rect 25340 14028 25396 14084
rect 25452 13970 25508 13972
rect 25452 13918 25454 13970
rect 25454 13918 25506 13970
rect 25506 13918 25508 13970
rect 25452 13916 25508 13918
rect 25228 13132 25284 13188
rect 23212 12348 23268 12404
rect 24332 11900 24388 11956
rect 24444 11788 24500 11844
rect 25228 11954 25284 11956
rect 25228 11902 25230 11954
rect 25230 11902 25282 11954
rect 25282 11902 25284 11954
rect 25228 11900 25284 11902
rect 25564 11954 25620 11956
rect 25564 11902 25566 11954
rect 25566 11902 25618 11954
rect 25618 11902 25620 11954
rect 25564 11900 25620 11902
rect 25004 11394 25060 11396
rect 25004 11342 25006 11394
rect 25006 11342 25058 11394
rect 25058 11342 25060 11394
rect 25004 11340 25060 11342
rect 21532 9884 21588 9940
rect 21868 10108 21924 10164
rect 21308 9714 21364 9716
rect 21308 9662 21310 9714
rect 21310 9662 21362 9714
rect 21362 9662 21364 9714
rect 21308 9660 21364 9662
rect 19852 8428 19908 8484
rect 23660 10108 23716 10164
rect 22204 9826 22260 9828
rect 22204 9774 22206 9826
rect 22206 9774 22258 9826
rect 22258 9774 22260 9826
rect 22204 9772 22260 9774
rect 23436 9884 23492 9940
rect 19404 7980 19460 8036
rect 20300 8370 20356 8372
rect 20300 8318 20302 8370
rect 20302 8318 20354 8370
rect 20354 8318 20356 8370
rect 20300 8316 20356 8318
rect 20524 8258 20580 8260
rect 20524 8206 20526 8258
rect 20526 8206 20578 8258
rect 20578 8206 20580 8258
rect 20524 8204 20580 8206
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 21308 8204 21364 8260
rect 21532 8146 21588 8148
rect 21532 8094 21534 8146
rect 21534 8094 21586 8146
rect 21586 8094 21588 8146
rect 21532 8092 21588 8094
rect 21420 7980 21476 8036
rect 21644 7756 21700 7812
rect 21532 6690 21588 6692
rect 21532 6638 21534 6690
rect 21534 6638 21586 6690
rect 21586 6638 21588 6690
rect 21532 6636 21588 6638
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 1708 5404 1764 5460
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 23660 9938 23716 9940
rect 23660 9886 23662 9938
rect 23662 9886 23714 9938
rect 23714 9886 23716 9938
rect 23660 9884 23716 9886
rect 22204 9324 22260 9380
rect 22092 8258 22148 8260
rect 22092 8206 22094 8258
rect 22094 8206 22146 8258
rect 22146 8206 22148 8258
rect 22092 8204 22148 8206
rect 21980 7756 22036 7812
rect 21868 6524 21924 6580
rect 21980 6636 22036 6692
rect 22764 9548 22820 9604
rect 22540 9212 22596 9268
rect 22428 7756 22484 7812
rect 21644 5292 21700 5348
rect 18844 5068 18900 5124
rect 19516 5068 19572 5124
rect 1708 4898 1764 4900
rect 1708 4846 1710 4898
rect 1710 4846 1762 4898
rect 1762 4846 1764 4898
rect 1708 4844 1764 4846
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19852 4508 19908 4564
rect 1708 4060 1764 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19516 3612 19572 3668
rect 1708 3388 1764 3444
rect 19628 3442 19684 3444
rect 19628 3390 19630 3442
rect 19630 3390 19682 3442
rect 19682 3390 19684 3442
rect 19628 3388 19684 3390
rect 22876 9324 22932 9380
rect 23772 9212 23828 9268
rect 23884 9154 23940 9156
rect 23884 9102 23886 9154
rect 23886 9102 23938 9154
rect 23938 9102 23940 9154
rect 23884 9100 23940 9102
rect 22764 8146 22820 8148
rect 22764 8094 22766 8146
rect 22766 8094 22818 8146
rect 22818 8094 22820 8146
rect 22764 8092 22820 8094
rect 24556 10556 24612 10612
rect 24444 9602 24500 9604
rect 24444 9550 24446 9602
rect 24446 9550 24498 9602
rect 24498 9550 24500 9602
rect 24444 9548 24500 9550
rect 24332 9436 24388 9492
rect 25900 14252 25956 14308
rect 25340 10610 25396 10612
rect 25340 10558 25342 10610
rect 25342 10558 25394 10610
rect 25394 10558 25396 10610
rect 25340 10556 25396 10558
rect 24780 9714 24836 9716
rect 24780 9662 24782 9714
rect 24782 9662 24834 9714
rect 24834 9662 24836 9714
rect 24780 9660 24836 9662
rect 24668 9212 24724 9268
rect 25564 9884 25620 9940
rect 25228 9602 25284 9604
rect 25228 9550 25230 9602
rect 25230 9550 25282 9602
rect 25282 9550 25284 9602
rect 25228 9548 25284 9550
rect 25676 9266 25732 9268
rect 25676 9214 25678 9266
rect 25678 9214 25730 9266
rect 25730 9214 25732 9266
rect 25676 9212 25732 9214
rect 25452 9154 25508 9156
rect 25452 9102 25454 9154
rect 25454 9102 25506 9154
rect 25506 9102 25508 9154
rect 25452 9100 25508 9102
rect 24668 9042 24724 9044
rect 24668 8990 24670 9042
rect 24670 8990 24722 9042
rect 24722 8990 24724 9042
rect 24668 8988 24724 8990
rect 24220 8092 24276 8148
rect 26012 13468 26068 13524
rect 26348 11900 26404 11956
rect 25900 9772 25956 9828
rect 26236 9996 26292 10052
rect 26348 9884 26404 9940
rect 26236 9324 26292 9380
rect 26348 9042 26404 9044
rect 26348 8990 26350 9042
rect 26350 8990 26402 9042
rect 26402 8990 26404 9042
rect 26348 8988 26404 8990
rect 26348 7980 26404 8036
rect 22540 6636 22596 6692
rect 22988 6578 23044 6580
rect 22988 6526 22990 6578
rect 22990 6526 23042 6578
rect 23042 6526 23044 6578
rect 22988 6524 23044 6526
rect 24108 6412 24164 6468
rect 23212 6130 23268 6132
rect 23212 6078 23214 6130
rect 23214 6078 23266 6130
rect 23266 6078 23268 6130
rect 23212 6076 23268 6078
rect 23436 6018 23492 6020
rect 23436 5966 23438 6018
rect 23438 5966 23490 6018
rect 23490 5966 23492 6018
rect 23436 5964 23492 5966
rect 24332 6578 24388 6580
rect 24332 6526 24334 6578
rect 24334 6526 24386 6578
rect 24386 6526 24388 6578
rect 24332 6524 24388 6526
rect 24220 5964 24276 6020
rect 23100 5292 23156 5348
rect 22876 5122 22932 5124
rect 22876 5070 22878 5122
rect 22878 5070 22930 5122
rect 22930 5070 22932 5122
rect 22876 5068 22932 5070
rect 24108 5068 24164 5124
rect 24892 6578 24948 6580
rect 24892 6526 24894 6578
rect 24894 6526 24946 6578
rect 24946 6526 24948 6578
rect 24892 6524 24948 6526
rect 25452 7644 25508 7700
rect 25452 6748 25508 6804
rect 25900 6300 25956 6356
rect 26012 6076 26068 6132
rect 25564 5906 25620 5908
rect 25564 5854 25566 5906
rect 25566 5854 25618 5906
rect 25618 5854 25620 5906
rect 25564 5852 25620 5854
rect 28140 20748 28196 20804
rect 27020 19964 27076 20020
rect 27244 20018 27300 20020
rect 27244 19966 27246 20018
rect 27246 19966 27298 20018
rect 27298 19966 27300 20018
rect 27244 19964 27300 19966
rect 27468 19906 27524 19908
rect 27468 19854 27470 19906
rect 27470 19854 27522 19906
rect 27522 19854 27524 19906
rect 27468 19852 27524 19854
rect 27020 19628 27076 19684
rect 27244 18450 27300 18452
rect 27244 18398 27246 18450
rect 27246 18398 27298 18450
rect 27298 18398 27300 18450
rect 27244 18396 27300 18398
rect 28476 22258 28532 22260
rect 28476 22206 28478 22258
rect 28478 22206 28530 22258
rect 28530 22206 28532 22258
rect 28476 22204 28532 22206
rect 29484 26850 29540 26852
rect 29484 26798 29486 26850
rect 29486 26798 29538 26850
rect 29538 26798 29540 26850
rect 29484 26796 29540 26798
rect 29932 26908 29988 26964
rect 29148 23212 29204 23268
rect 29036 22594 29092 22596
rect 29036 22542 29038 22594
rect 29038 22542 29090 22594
rect 29090 22542 29092 22594
rect 29036 22540 29092 22542
rect 31388 32172 31444 32228
rect 31612 32620 31668 32676
rect 31500 32508 31556 32564
rect 32172 37826 32228 37828
rect 32172 37774 32174 37826
rect 32174 37774 32226 37826
rect 32226 37774 32228 37826
rect 32172 37772 32228 37774
rect 31836 35756 31892 35812
rect 32060 37378 32116 37380
rect 32060 37326 32062 37378
rect 32062 37326 32114 37378
rect 32114 37326 32116 37378
rect 32060 37324 32116 37326
rect 32508 37826 32564 37828
rect 32508 37774 32510 37826
rect 32510 37774 32562 37826
rect 32562 37774 32564 37826
rect 32508 37772 32564 37774
rect 32508 37212 32564 37268
rect 32396 36988 32452 37044
rect 32284 35810 32340 35812
rect 32284 35758 32286 35810
rect 32286 35758 32338 35810
rect 32338 35758 32340 35810
rect 32284 35756 32340 35758
rect 32508 35698 32564 35700
rect 32508 35646 32510 35698
rect 32510 35646 32562 35698
rect 32562 35646 32564 35698
rect 32508 35644 32564 35646
rect 32172 35420 32228 35476
rect 32396 34300 32452 34356
rect 32284 34130 32340 34132
rect 32284 34078 32286 34130
rect 32286 34078 32338 34130
rect 32338 34078 32340 34130
rect 32284 34076 32340 34078
rect 32172 33570 32228 33572
rect 32172 33518 32174 33570
rect 32174 33518 32226 33570
rect 32226 33518 32228 33570
rect 32172 33516 32228 33518
rect 32284 33404 32340 33460
rect 31836 32844 31892 32900
rect 32172 32732 32228 32788
rect 31836 31724 31892 31780
rect 32060 30322 32116 30324
rect 32060 30270 32062 30322
rect 32062 30270 32114 30322
rect 32114 30270 32116 30322
rect 32060 30268 32116 30270
rect 32172 30156 32228 30212
rect 30828 29426 30884 29428
rect 30828 29374 30830 29426
rect 30830 29374 30882 29426
rect 30882 29374 30884 29426
rect 30828 29372 30884 29374
rect 30940 28700 30996 28756
rect 31836 29820 31892 29876
rect 31948 29708 32004 29764
rect 31500 29372 31556 29428
rect 31276 28642 31332 28644
rect 31276 28590 31278 28642
rect 31278 28590 31330 28642
rect 31330 28590 31332 28642
rect 31276 28588 31332 28590
rect 40348 39004 40404 39060
rect 33180 38722 33236 38724
rect 33180 38670 33182 38722
rect 33182 38670 33234 38722
rect 33234 38670 33236 38722
rect 33180 38668 33236 38670
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 40124 38332 40180 38388
rect 33292 37772 33348 37828
rect 40124 37660 40180 37716
rect 32732 30156 32788 30212
rect 32844 36988 32900 37044
rect 32396 29596 32452 29652
rect 40124 36988 40180 37044
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 33068 35698 33124 35700
rect 33068 35646 33070 35698
rect 33070 35646 33122 35698
rect 33122 35646 33124 35698
rect 33068 35644 33124 35646
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 33516 33292 33572 33348
rect 33404 32396 33460 32452
rect 33964 32450 34020 32452
rect 33964 32398 33966 32450
rect 33966 32398 34018 32450
rect 34018 32398 34020 32450
rect 33964 32396 34020 32398
rect 33628 32284 33684 32340
rect 32956 30210 33012 30212
rect 32956 30158 32958 30210
rect 32958 30158 33010 30210
rect 33010 30158 33012 30210
rect 32956 30156 33012 30158
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34412 33292 34468 33348
rect 34972 33234 35028 33236
rect 34972 33182 34974 33234
rect 34974 33182 35026 33234
rect 35026 33182 35028 33234
rect 34972 33180 35028 33182
rect 35868 33234 35924 33236
rect 35868 33182 35870 33234
rect 35870 33182 35922 33234
rect 35922 33182 35924 33234
rect 35868 33180 35924 33182
rect 35756 33122 35812 33124
rect 35756 33070 35758 33122
rect 35758 33070 35810 33122
rect 35810 33070 35812 33122
rect 35756 33068 35812 33070
rect 33964 30210 34020 30212
rect 33964 30158 33966 30210
rect 33966 30158 34018 30210
rect 34018 30158 34020 30210
rect 33964 30156 34020 30158
rect 34188 32284 34244 32340
rect 34188 31276 34244 31332
rect 32844 29820 32900 29876
rect 33292 29708 33348 29764
rect 32172 28588 32228 28644
rect 31164 27356 31220 27412
rect 31612 27186 31668 27188
rect 31612 27134 31614 27186
rect 31614 27134 31666 27186
rect 31666 27134 31668 27186
rect 31612 27132 31668 27134
rect 31388 26962 31444 26964
rect 31388 26910 31390 26962
rect 31390 26910 31442 26962
rect 31442 26910 31444 26962
rect 31388 26908 31444 26910
rect 32284 27970 32340 27972
rect 32284 27918 32286 27970
rect 32286 27918 32338 27970
rect 32338 27918 32340 27970
rect 32284 27916 32340 27918
rect 31724 27020 31780 27076
rect 30940 26290 30996 26292
rect 30940 26238 30942 26290
rect 30942 26238 30994 26290
rect 30994 26238 30996 26290
rect 30940 26236 30996 26238
rect 31500 26066 31556 26068
rect 31500 26014 31502 26066
rect 31502 26014 31554 26066
rect 31554 26014 31556 26066
rect 31500 26012 31556 26014
rect 31164 25618 31220 25620
rect 31164 25566 31166 25618
rect 31166 25566 31218 25618
rect 31218 25566 31220 25618
rect 31164 25564 31220 25566
rect 30268 25506 30324 25508
rect 30268 25454 30270 25506
rect 30270 25454 30322 25506
rect 30322 25454 30324 25506
rect 30268 25452 30324 25454
rect 30828 25452 30884 25508
rect 30492 23324 30548 23380
rect 30044 23266 30100 23268
rect 30044 23214 30046 23266
rect 30046 23214 30098 23266
rect 30098 23214 30100 23266
rect 30044 23212 30100 23214
rect 29932 23042 29988 23044
rect 29932 22990 29934 23042
rect 29934 22990 29986 23042
rect 29986 22990 29988 23042
rect 29932 22988 29988 22990
rect 29148 22146 29204 22148
rect 29148 22094 29150 22146
rect 29150 22094 29202 22146
rect 29202 22094 29204 22146
rect 29148 22092 29204 22094
rect 28812 21586 28868 21588
rect 28812 21534 28814 21586
rect 28814 21534 28866 21586
rect 28866 21534 28868 21586
rect 28812 21532 28868 21534
rect 28364 19964 28420 20020
rect 28140 19740 28196 19796
rect 28700 19516 28756 19572
rect 28588 19234 28644 19236
rect 28588 19182 28590 19234
rect 28590 19182 28642 19234
rect 28642 19182 28644 19234
rect 28588 19180 28644 19182
rect 27132 17554 27188 17556
rect 27132 17502 27134 17554
rect 27134 17502 27186 17554
rect 27186 17502 27188 17554
rect 27132 17500 27188 17502
rect 27916 16268 27972 16324
rect 27244 14588 27300 14644
rect 26796 14252 26852 14308
rect 27132 14476 27188 14532
rect 26684 13580 26740 13636
rect 27468 13468 27524 13524
rect 27244 13186 27300 13188
rect 27244 13134 27246 13186
rect 27246 13134 27298 13186
rect 27298 13134 27300 13186
rect 27244 13132 27300 13134
rect 26908 9212 26964 9268
rect 27132 9324 27188 9380
rect 28476 16940 28532 16996
rect 28588 16268 28644 16324
rect 28700 14812 28756 14868
rect 28812 13916 28868 13972
rect 28252 13580 28308 13636
rect 29260 19404 29316 19460
rect 29596 21698 29652 21700
rect 29596 21646 29598 21698
rect 29598 21646 29650 21698
rect 29650 21646 29652 21698
rect 29596 21644 29652 21646
rect 29596 21362 29652 21364
rect 29596 21310 29598 21362
rect 29598 21310 29650 21362
rect 29650 21310 29652 21362
rect 29596 21308 29652 21310
rect 29932 22092 29988 22148
rect 29484 20802 29540 20804
rect 29484 20750 29486 20802
rect 29486 20750 29538 20802
rect 29538 20750 29540 20802
rect 29484 20748 29540 20750
rect 29372 20076 29428 20132
rect 29820 20972 29876 21028
rect 30828 21026 30884 21028
rect 30828 20974 30830 21026
rect 30830 20974 30882 21026
rect 30882 20974 30884 21026
rect 30828 20972 30884 20974
rect 29932 20018 29988 20020
rect 29932 19966 29934 20018
rect 29934 19966 29986 20018
rect 29986 19966 29988 20018
rect 29932 19964 29988 19966
rect 30380 19964 30436 20020
rect 29484 19516 29540 19572
rect 29260 19180 29316 19236
rect 29148 17666 29204 17668
rect 29148 17614 29150 17666
rect 29150 17614 29202 17666
rect 29202 17614 29204 17666
rect 29148 17612 29204 17614
rect 29148 16994 29204 16996
rect 29148 16942 29150 16994
rect 29150 16942 29202 16994
rect 29202 16942 29204 16994
rect 29148 16940 29204 16942
rect 30604 19122 30660 19124
rect 30604 19070 30606 19122
rect 30606 19070 30658 19122
rect 30658 19070 30660 19122
rect 30604 19068 30660 19070
rect 29820 18620 29876 18676
rect 29484 17612 29540 17668
rect 30492 17554 30548 17556
rect 30492 17502 30494 17554
rect 30494 17502 30546 17554
rect 30546 17502 30548 17554
rect 30492 17500 30548 17502
rect 30716 17388 30772 17444
rect 29932 16940 29988 16996
rect 30156 16156 30212 16212
rect 29484 15820 29540 15876
rect 30044 15148 30100 15204
rect 29932 15036 29988 15092
rect 30156 15036 30212 15092
rect 29820 14700 29876 14756
rect 29148 14642 29204 14644
rect 29148 14590 29150 14642
rect 29150 14590 29202 14642
rect 29202 14590 29204 14642
rect 29148 14588 29204 14590
rect 29820 13970 29876 13972
rect 29820 13918 29822 13970
rect 29822 13918 29874 13970
rect 29874 13918 29876 13970
rect 29820 13916 29876 13918
rect 28924 13244 28980 13300
rect 27916 13132 27972 13188
rect 28028 12178 28084 12180
rect 28028 12126 28030 12178
rect 28030 12126 28082 12178
rect 28082 12126 28084 12178
rect 28028 12124 28084 12126
rect 28588 12178 28644 12180
rect 28588 12126 28590 12178
rect 28590 12126 28642 12178
rect 28642 12126 28644 12178
rect 28588 12124 28644 12126
rect 30156 13916 30212 13972
rect 30492 16994 30548 16996
rect 30492 16942 30494 16994
rect 30494 16942 30546 16994
rect 30546 16942 30548 16994
rect 30492 16940 30548 16942
rect 30828 16044 30884 16100
rect 30380 13804 30436 13860
rect 30492 14812 30548 14868
rect 31612 25394 31668 25396
rect 31612 25342 31614 25394
rect 31614 25342 31666 25394
rect 31666 25342 31668 25394
rect 31612 25340 31668 25342
rect 32060 27858 32116 27860
rect 32060 27806 32062 27858
rect 32062 27806 32114 27858
rect 32114 27806 32116 27858
rect 32060 27804 32116 27806
rect 33628 29372 33684 29428
rect 34076 29820 34132 29876
rect 33852 29148 33908 29204
rect 33068 28082 33124 28084
rect 33068 28030 33070 28082
rect 33070 28030 33122 28082
rect 33122 28030 33124 28082
rect 33068 28028 33124 28030
rect 31948 27634 32004 27636
rect 31948 27582 31950 27634
rect 31950 27582 32002 27634
rect 32002 27582 32004 27634
rect 31948 27580 32004 27582
rect 32060 27468 32116 27524
rect 32284 27356 32340 27412
rect 33516 27244 33572 27300
rect 33852 27804 33908 27860
rect 33068 26962 33124 26964
rect 33068 26910 33070 26962
rect 33070 26910 33122 26962
rect 33122 26910 33124 26962
rect 33068 26908 33124 26910
rect 32060 26290 32116 26292
rect 32060 26238 32062 26290
rect 32062 26238 32114 26290
rect 32114 26238 32116 26290
rect 32060 26236 32116 26238
rect 31388 24722 31444 24724
rect 31388 24670 31390 24722
rect 31390 24670 31442 24722
rect 31442 24670 31444 24722
rect 31388 24668 31444 24670
rect 32620 26460 32676 26516
rect 32844 26796 32900 26852
rect 32732 26012 32788 26068
rect 32172 25340 32228 25396
rect 32060 23548 32116 23604
rect 31276 22428 31332 22484
rect 31724 21644 31780 21700
rect 32172 21532 32228 21588
rect 31388 19964 31444 20020
rect 31836 20524 31892 20580
rect 31724 19740 31780 19796
rect 32508 20748 32564 20804
rect 32956 25116 33012 25172
rect 33740 26908 33796 26964
rect 33292 26514 33348 26516
rect 33292 26462 33294 26514
rect 33294 26462 33346 26514
rect 33346 26462 33348 26514
rect 33292 26460 33348 26462
rect 33292 26290 33348 26292
rect 33292 26238 33294 26290
rect 33294 26238 33346 26290
rect 33346 26238 33348 26290
rect 33292 26236 33348 26238
rect 33292 25116 33348 25172
rect 32956 24722 33012 24724
rect 32956 24670 32958 24722
rect 32958 24670 33010 24722
rect 33010 24670 33012 24722
rect 32956 24668 33012 24670
rect 33852 25340 33908 25396
rect 34076 23996 34132 24052
rect 33740 23548 33796 23604
rect 33740 23212 33796 23268
rect 32732 21532 32788 21588
rect 32620 20636 32676 20692
rect 31276 19516 31332 19572
rect 31276 19122 31332 19124
rect 31276 19070 31278 19122
rect 31278 19070 31330 19122
rect 31330 19070 31332 19122
rect 31276 19068 31332 19070
rect 31500 17612 31556 17668
rect 31164 17554 31220 17556
rect 31164 17502 31166 17554
rect 31166 17502 31218 17554
rect 31218 17502 31220 17554
rect 31164 17500 31220 17502
rect 32508 20018 32564 20020
rect 32508 19966 32510 20018
rect 32510 19966 32562 20018
rect 32562 19966 32564 20018
rect 32508 19964 32564 19966
rect 33404 22482 33460 22484
rect 33404 22430 33406 22482
rect 33406 22430 33458 22482
rect 33458 22430 33460 22482
rect 33404 22428 33460 22430
rect 33292 22316 33348 22372
rect 33068 22258 33124 22260
rect 33068 22206 33070 22258
rect 33070 22206 33122 22258
rect 33122 22206 33124 22258
rect 33068 22204 33124 22206
rect 33404 22092 33460 22148
rect 33516 21980 33572 22036
rect 33180 21586 33236 21588
rect 33180 21534 33182 21586
rect 33182 21534 33234 21586
rect 33234 21534 33236 21586
rect 33180 21532 33236 21534
rect 34636 31890 34692 31892
rect 34636 31838 34638 31890
rect 34638 31838 34690 31890
rect 34690 31838 34692 31890
rect 34636 31836 34692 31838
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35308 31500 35364 31556
rect 35644 32450 35700 32452
rect 35644 32398 35646 32450
rect 35646 32398 35698 32450
rect 35698 32398 35700 32450
rect 35644 32396 35700 32398
rect 35756 31778 35812 31780
rect 35756 31726 35758 31778
rect 35758 31726 35810 31778
rect 35810 31726 35812 31778
rect 35756 31724 35812 31726
rect 35980 31724 36036 31780
rect 35868 31218 35924 31220
rect 35868 31166 35870 31218
rect 35870 31166 35922 31218
rect 35922 31166 35924 31218
rect 35868 31164 35924 31166
rect 35084 31106 35140 31108
rect 35084 31054 35086 31106
rect 35086 31054 35138 31106
rect 35138 31054 35140 31106
rect 35084 31052 35140 31054
rect 35644 30882 35700 30884
rect 35644 30830 35646 30882
rect 35646 30830 35698 30882
rect 35698 30830 35700 30882
rect 35644 30828 35700 30830
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34636 30322 34692 30324
rect 34636 30270 34638 30322
rect 34638 30270 34690 30322
rect 34690 30270 34692 30322
rect 34636 30268 34692 30270
rect 35868 30268 35924 30324
rect 34524 30098 34580 30100
rect 34524 30046 34526 30098
rect 34526 30046 34578 30098
rect 34578 30046 34580 30098
rect 34524 30044 34580 30046
rect 35532 29148 35588 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35644 29372 35700 29428
rect 34412 28364 34468 28420
rect 35532 28418 35588 28420
rect 35532 28366 35534 28418
rect 35534 28366 35586 28418
rect 35586 28366 35588 28418
rect 35532 28364 35588 28366
rect 35420 27580 35476 27636
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35308 27298 35364 27300
rect 35308 27246 35310 27298
rect 35310 27246 35362 27298
rect 35362 27246 35364 27298
rect 35308 27244 35364 27246
rect 34860 27186 34916 27188
rect 34860 27134 34862 27186
rect 34862 27134 34914 27186
rect 34914 27134 34916 27186
rect 34860 27132 34916 27134
rect 34748 27020 34804 27076
rect 34524 26962 34580 26964
rect 34524 26910 34526 26962
rect 34526 26910 34578 26962
rect 34578 26910 34580 26962
rect 34524 26908 34580 26910
rect 35420 27074 35476 27076
rect 35420 27022 35422 27074
rect 35422 27022 35474 27074
rect 35474 27022 35476 27074
rect 35420 27020 35476 27022
rect 35308 26178 35364 26180
rect 35308 26126 35310 26178
rect 35310 26126 35362 26178
rect 35362 26126 35364 26178
rect 35308 26124 35364 26126
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 36652 32562 36708 32564
rect 36652 32510 36654 32562
rect 36654 32510 36706 32562
rect 36706 32510 36708 32562
rect 36652 32508 36708 32510
rect 37772 33068 37828 33124
rect 37100 32508 37156 32564
rect 36428 31948 36484 32004
rect 36764 31836 36820 31892
rect 36316 31500 36372 31556
rect 36540 31612 36596 31668
rect 36316 31276 36372 31332
rect 36204 30156 36260 30212
rect 35980 29986 36036 29988
rect 35980 29934 35982 29986
rect 35982 29934 36034 29986
rect 36034 29934 36036 29986
rect 35980 29932 36036 29934
rect 36876 31948 36932 32004
rect 36988 31836 37044 31892
rect 37884 31890 37940 31892
rect 37884 31838 37886 31890
rect 37886 31838 37938 31890
rect 37938 31838 37940 31890
rect 37884 31836 37940 31838
rect 37100 31778 37156 31780
rect 37100 31726 37102 31778
rect 37102 31726 37154 31778
rect 37154 31726 37156 31778
rect 37100 31724 37156 31726
rect 37548 31666 37604 31668
rect 37548 31614 37550 31666
rect 37550 31614 37602 31666
rect 37602 31614 37604 31666
rect 37548 31612 37604 31614
rect 37212 31500 37268 31556
rect 36876 29932 36932 29988
rect 35868 29426 35924 29428
rect 35868 29374 35870 29426
rect 35870 29374 35922 29426
rect 35922 29374 35924 29426
rect 35868 29372 35924 29374
rect 36316 27244 36372 27300
rect 36316 26796 36372 26852
rect 34188 23324 34244 23380
rect 34188 22316 34244 22372
rect 34412 22258 34468 22260
rect 34412 22206 34414 22258
rect 34414 22206 34466 22258
rect 34466 22206 34468 22258
rect 34412 22204 34468 22206
rect 33852 21532 33908 21588
rect 33292 21420 33348 21476
rect 34188 21474 34244 21476
rect 34188 21422 34190 21474
rect 34190 21422 34242 21474
rect 34242 21422 34244 21474
rect 34188 21420 34244 21422
rect 33292 20524 33348 20580
rect 33404 20076 33460 20132
rect 32956 19964 33012 20020
rect 33516 20018 33572 20020
rect 33516 19966 33518 20018
rect 33518 19966 33570 20018
rect 33570 19966 33572 20018
rect 33516 19964 33572 19966
rect 32956 19122 33012 19124
rect 32956 19070 32958 19122
rect 32958 19070 33010 19122
rect 33010 19070 33012 19122
rect 32956 19068 33012 19070
rect 34188 20802 34244 20804
rect 34188 20750 34190 20802
rect 34190 20750 34242 20802
rect 34242 20750 34244 20802
rect 34188 20748 34244 20750
rect 34636 22146 34692 22148
rect 34636 22094 34638 22146
rect 34638 22094 34690 22146
rect 34690 22094 34692 22146
rect 34636 22092 34692 22094
rect 34860 21698 34916 21700
rect 34860 21646 34862 21698
rect 34862 21646 34914 21698
rect 34914 21646 34916 21698
rect 34860 21644 34916 21646
rect 34748 20690 34804 20692
rect 34748 20638 34750 20690
rect 34750 20638 34802 20690
rect 34802 20638 34804 20690
rect 34748 20636 34804 20638
rect 34524 20524 34580 20580
rect 33852 20300 33908 20356
rect 34188 20300 34244 20356
rect 33740 20018 33796 20020
rect 33740 19966 33742 20018
rect 33742 19966 33794 20018
rect 33794 19966 33796 20018
rect 33740 19964 33796 19966
rect 33628 18844 33684 18900
rect 33852 19740 33908 19796
rect 34860 20018 34916 20020
rect 34860 19966 34862 20018
rect 34862 19966 34914 20018
rect 34914 19966 34916 20018
rect 34860 19964 34916 19966
rect 37660 30828 37716 30884
rect 37324 30210 37380 30212
rect 37324 30158 37326 30210
rect 37326 30158 37378 30210
rect 37378 30158 37380 30210
rect 37324 30156 37380 30158
rect 37884 29986 37940 29988
rect 37884 29934 37886 29986
rect 37886 29934 37938 29986
rect 37938 29934 37940 29986
rect 37884 29932 37940 29934
rect 37884 29484 37940 29540
rect 40124 30268 40180 30324
rect 38444 29986 38500 29988
rect 38444 29934 38446 29986
rect 38446 29934 38498 29986
rect 38498 29934 38500 29986
rect 38444 29932 38500 29934
rect 38220 29372 38276 29428
rect 35756 24556 35812 24612
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 38556 29260 38612 29316
rect 40124 29314 40180 29316
rect 40124 29262 40126 29314
rect 40126 29262 40178 29314
rect 40178 29262 40180 29314
rect 40124 29260 40180 29262
rect 37996 27298 38052 27300
rect 37996 27246 37998 27298
rect 37998 27246 38050 27298
rect 38050 27246 38052 27298
rect 37996 27244 38052 27246
rect 36764 23996 36820 24052
rect 36540 23938 36596 23940
rect 36540 23886 36542 23938
rect 36542 23886 36594 23938
rect 36594 23886 36596 23938
rect 36540 23884 36596 23886
rect 37212 23938 37268 23940
rect 37212 23886 37214 23938
rect 37214 23886 37266 23938
rect 37266 23886 37268 23938
rect 37212 23884 37268 23886
rect 36652 23378 36708 23380
rect 36652 23326 36654 23378
rect 36654 23326 36706 23378
rect 36706 23326 36708 23378
rect 36652 23324 36708 23326
rect 35084 21644 35140 21700
rect 35532 22316 35588 22372
rect 35868 22204 35924 22260
rect 35196 21980 35252 22036
rect 35532 21644 35588 21700
rect 35420 21586 35476 21588
rect 35420 21534 35422 21586
rect 35422 21534 35474 21586
rect 35474 21534 35476 21586
rect 35420 21532 35476 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 32508 18396 32564 18452
rect 33740 18508 33796 18564
rect 34076 18172 34132 18228
rect 34412 19068 34468 19124
rect 34300 18396 34356 18452
rect 32172 17442 32228 17444
rect 32172 17390 32174 17442
rect 32174 17390 32226 17442
rect 32226 17390 32228 17442
rect 32172 17388 32228 17390
rect 31948 16940 32004 16996
rect 32844 16716 32900 16772
rect 31948 15986 32004 15988
rect 31948 15934 31950 15986
rect 31950 15934 32002 15986
rect 32002 15934 32004 15986
rect 31948 15932 32004 15934
rect 31052 15260 31108 15316
rect 31052 15090 31108 15092
rect 31052 15038 31054 15090
rect 31054 15038 31106 15090
rect 31106 15038 31108 15090
rect 31052 15036 31108 15038
rect 31164 14924 31220 14980
rect 30940 14812 30996 14868
rect 30604 13356 30660 13412
rect 30716 13468 30772 13524
rect 31388 15314 31444 15316
rect 31388 15262 31390 15314
rect 31390 15262 31442 15314
rect 31442 15262 31444 15314
rect 31388 15260 31444 15262
rect 31612 14924 31668 14980
rect 32844 15484 32900 15540
rect 33068 17500 33124 17556
rect 33852 17554 33908 17556
rect 33852 17502 33854 17554
rect 33854 17502 33906 17554
rect 33906 17502 33908 17554
rect 33852 17500 33908 17502
rect 33404 17106 33460 17108
rect 33404 17054 33406 17106
rect 33406 17054 33458 17106
rect 33458 17054 33460 17106
rect 33404 17052 33460 17054
rect 33852 17052 33908 17108
rect 33516 16716 33572 16772
rect 33068 15932 33124 15988
rect 33292 15596 33348 15652
rect 32172 15314 32228 15316
rect 32172 15262 32174 15314
rect 32174 15262 32226 15314
rect 32226 15262 32228 15314
rect 32172 15260 32228 15262
rect 32060 14700 32116 14756
rect 32172 14028 32228 14084
rect 31612 13468 31668 13524
rect 31388 13356 31444 13412
rect 31052 12962 31108 12964
rect 31052 12910 31054 12962
rect 31054 12910 31106 12962
rect 31106 12910 31108 12962
rect 31052 12908 31108 12910
rect 31164 12796 31220 12852
rect 29820 12124 29876 12180
rect 28252 11282 28308 11284
rect 28252 11230 28254 11282
rect 28254 11230 28306 11282
rect 28306 11230 28308 11282
rect 28252 11228 28308 11230
rect 27916 11170 27972 11172
rect 27916 11118 27918 11170
rect 27918 11118 27970 11170
rect 27970 11118 27972 11170
rect 27916 11116 27972 11118
rect 28588 11116 28644 11172
rect 28252 10668 28308 10724
rect 27692 9100 27748 9156
rect 28140 9266 28196 9268
rect 28140 9214 28142 9266
rect 28142 9214 28194 9266
rect 28194 9214 28196 9266
rect 28140 9212 28196 9214
rect 28924 10722 28980 10724
rect 28924 10670 28926 10722
rect 28926 10670 28978 10722
rect 28978 10670 28980 10722
rect 28924 10668 28980 10670
rect 29484 11282 29540 11284
rect 29484 11230 29486 11282
rect 29486 11230 29538 11282
rect 29538 11230 29540 11282
rect 29484 11228 29540 11230
rect 30044 11228 30100 11284
rect 29708 10668 29764 10724
rect 29484 10556 29540 10612
rect 32060 13580 32116 13636
rect 30940 11340 30996 11396
rect 30828 11116 30884 11172
rect 30268 10610 30324 10612
rect 30268 10558 30270 10610
rect 30270 10558 30322 10610
rect 30322 10558 30324 10610
rect 30268 10556 30324 10558
rect 29148 9266 29204 9268
rect 29148 9214 29150 9266
rect 29150 9214 29202 9266
rect 29202 9214 29204 9266
rect 29148 9212 29204 9214
rect 26460 6748 26516 6804
rect 28252 8428 28308 8484
rect 27580 7980 27636 8036
rect 28364 8034 28420 8036
rect 28364 7982 28366 8034
rect 28366 7982 28418 8034
rect 28418 7982 28420 8034
rect 28364 7980 28420 7982
rect 27468 6860 27524 6916
rect 28364 6860 28420 6916
rect 27132 6466 27188 6468
rect 27132 6414 27134 6466
rect 27134 6414 27186 6466
rect 27186 6414 27188 6466
rect 27132 6412 27188 6414
rect 26348 6300 26404 6356
rect 31612 12178 31668 12180
rect 31612 12126 31614 12178
rect 31614 12126 31666 12178
rect 31666 12126 31668 12178
rect 31612 12124 31668 12126
rect 32172 13132 32228 13188
rect 33068 13804 33124 13860
rect 32508 13356 32564 13412
rect 33068 13186 33124 13188
rect 33068 13134 33070 13186
rect 33070 13134 33122 13186
rect 33122 13134 33124 13186
rect 33068 13132 33124 13134
rect 32620 12962 32676 12964
rect 32620 12910 32622 12962
rect 32622 12910 32674 12962
rect 32674 12910 32676 12962
rect 32620 12908 32676 12910
rect 31724 11228 31780 11284
rect 31388 11116 31444 11172
rect 31836 11116 31892 11172
rect 29596 9548 29652 9604
rect 30380 9602 30436 9604
rect 30380 9550 30382 9602
rect 30382 9550 30434 9602
rect 30434 9550 30436 9602
rect 30380 9548 30436 9550
rect 31388 9772 31444 9828
rect 31724 10332 31780 10388
rect 30940 9212 30996 9268
rect 34188 16716 34244 16772
rect 34636 18562 34692 18564
rect 34636 18510 34638 18562
rect 34638 18510 34690 18562
rect 34690 18510 34692 18562
rect 34636 18508 34692 18510
rect 35420 20018 35476 20020
rect 35420 19966 35422 20018
rect 35422 19966 35474 20018
rect 35474 19966 35476 20018
rect 35420 19964 35476 19966
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34860 18338 34916 18340
rect 34860 18286 34862 18338
rect 34862 18286 34914 18338
rect 34914 18286 34916 18338
rect 34860 18284 34916 18286
rect 34636 18172 34692 18228
rect 34524 17890 34580 17892
rect 34524 17838 34526 17890
rect 34526 17838 34578 17890
rect 34578 17838 34580 17890
rect 34524 17836 34580 17838
rect 34300 17276 34356 17332
rect 34636 16940 34692 16996
rect 36092 21644 36148 21700
rect 37324 22370 37380 22372
rect 37324 22318 37326 22370
rect 37326 22318 37378 22370
rect 37378 22318 37380 22370
rect 37324 22316 37380 22318
rect 36316 22092 36372 22148
rect 36876 22092 36932 22148
rect 36428 21810 36484 21812
rect 36428 21758 36430 21810
rect 36430 21758 36482 21810
rect 36482 21758 36484 21810
rect 36428 21756 36484 21758
rect 36428 20188 36484 20244
rect 36988 21644 37044 21700
rect 37212 21644 37268 21700
rect 37212 20188 37268 20244
rect 36876 19964 36932 20020
rect 39564 26796 39620 26852
rect 39788 26572 39844 26628
rect 40124 26796 40180 26852
rect 40012 26236 40068 26292
rect 39788 25228 39844 25284
rect 40124 24610 40180 24612
rect 40124 24558 40126 24610
rect 40126 24558 40178 24610
rect 40178 24558 40180 24610
rect 40124 24556 40180 24558
rect 40124 24050 40180 24052
rect 40124 23998 40126 24050
rect 40126 23998 40178 24050
rect 40178 23998 40180 24050
rect 40124 23996 40180 23998
rect 38332 23324 38388 23380
rect 38444 22146 38500 22148
rect 38444 22094 38446 22146
rect 38446 22094 38498 22146
rect 38498 22094 38500 22146
rect 38444 22092 38500 22094
rect 38556 21644 38612 21700
rect 38108 21586 38164 21588
rect 38108 21534 38110 21586
rect 38110 21534 38162 21586
rect 38162 21534 38164 21586
rect 38108 21532 38164 21534
rect 37436 21362 37492 21364
rect 37436 21310 37438 21362
rect 37438 21310 37490 21362
rect 37490 21310 37492 21362
rect 37436 21308 37492 21310
rect 35308 18172 35364 18228
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34972 17052 35028 17108
rect 34748 16828 34804 16884
rect 35084 17388 35140 17444
rect 36540 19180 36596 19236
rect 38892 20130 38948 20132
rect 38892 20078 38894 20130
rect 38894 20078 38946 20130
rect 38946 20078 38948 20130
rect 38892 20076 38948 20078
rect 40124 21532 40180 21588
rect 40012 20860 40068 20916
rect 39676 20130 39732 20132
rect 39676 20078 39678 20130
rect 39678 20078 39730 20130
rect 39730 20078 39732 20130
rect 39676 20076 39732 20078
rect 39116 19740 39172 19796
rect 40012 19516 40068 19572
rect 37436 19234 37492 19236
rect 37436 19182 37438 19234
rect 37438 19182 37490 19234
rect 37490 19182 37492 19234
rect 37436 19180 37492 19182
rect 36652 18562 36708 18564
rect 36652 18510 36654 18562
rect 36654 18510 36706 18562
rect 36706 18510 36708 18562
rect 36652 18508 36708 18510
rect 37324 18674 37380 18676
rect 37324 18622 37326 18674
rect 37326 18622 37378 18674
rect 37378 18622 37380 18674
rect 37324 18620 37380 18622
rect 36988 18396 37044 18452
rect 36316 18338 36372 18340
rect 36316 18286 36318 18338
rect 36318 18286 36370 18338
rect 36370 18286 36372 18338
rect 36316 18284 36372 18286
rect 36092 17836 36148 17892
rect 35532 16882 35588 16884
rect 35532 16830 35534 16882
rect 35534 16830 35586 16882
rect 35586 16830 35588 16882
rect 35532 16828 35588 16830
rect 35980 17052 36036 17108
rect 35196 16770 35252 16772
rect 35196 16718 35198 16770
rect 35198 16718 35250 16770
rect 35250 16718 35252 16770
rect 35196 16716 35252 16718
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35084 16268 35140 16324
rect 34300 15596 34356 15652
rect 33404 14700 33460 14756
rect 33516 14028 33572 14084
rect 33292 13132 33348 13188
rect 33516 12124 33572 12180
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34636 13804 34692 13860
rect 35644 13858 35700 13860
rect 35644 13806 35646 13858
rect 35646 13806 35698 13858
rect 35698 13806 35700 13858
rect 35644 13804 35700 13806
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 33964 13132 34020 13188
rect 34076 12796 34132 12852
rect 35644 12850 35700 12852
rect 35644 12798 35646 12850
rect 35646 12798 35698 12850
rect 35698 12798 35700 12850
rect 35644 12796 35700 12798
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 32956 11394 33012 11396
rect 32956 11342 32958 11394
rect 32958 11342 33010 11394
rect 33010 11342 33012 11394
rect 32956 11340 33012 11342
rect 33516 11340 33572 11396
rect 32732 10332 32788 10388
rect 32844 11228 32900 11284
rect 33292 11282 33348 11284
rect 33292 11230 33294 11282
rect 33294 11230 33346 11282
rect 33346 11230 33348 11282
rect 33292 11228 33348 11230
rect 34076 10444 34132 10500
rect 32844 9938 32900 9940
rect 32844 9886 32846 9938
rect 32846 9886 32898 9938
rect 32898 9886 32900 9938
rect 32844 9884 32900 9886
rect 33852 9884 33908 9940
rect 35644 10498 35700 10500
rect 35644 10446 35646 10498
rect 35646 10446 35698 10498
rect 35698 10446 35700 10498
rect 35644 10444 35700 10446
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34188 9826 34244 9828
rect 34188 9774 34190 9826
rect 34190 9774 34242 9826
rect 34242 9774 34244 9826
rect 34188 9772 34244 9774
rect 34748 9772 34804 9828
rect 32284 9660 32340 9716
rect 31948 9602 32004 9604
rect 31948 9550 31950 9602
rect 31950 9550 32002 9602
rect 32002 9550 32004 9602
rect 31948 9548 32004 9550
rect 29596 8428 29652 8484
rect 33292 9714 33348 9716
rect 33292 9662 33294 9714
rect 33294 9662 33346 9714
rect 33346 9662 33348 9714
rect 33292 9660 33348 9662
rect 34524 9714 34580 9716
rect 34524 9662 34526 9714
rect 34526 9662 34578 9714
rect 34578 9662 34580 9714
rect 34524 9660 34580 9662
rect 32396 9548 32452 9604
rect 33068 9548 33124 9604
rect 32508 9042 32564 9044
rect 32508 8990 32510 9042
rect 32510 8990 32562 9042
rect 32562 8990 32564 9042
rect 32508 8988 32564 8990
rect 29372 6860 29428 6916
rect 37772 18508 37828 18564
rect 37436 18284 37492 18340
rect 36764 17106 36820 17108
rect 36764 17054 36766 17106
rect 36766 17054 36818 17106
rect 36818 17054 36820 17106
rect 36764 17052 36820 17054
rect 36652 16994 36708 16996
rect 36652 16942 36654 16994
rect 36654 16942 36706 16994
rect 36706 16942 36708 16994
rect 36652 16940 36708 16942
rect 36204 16828 36260 16884
rect 37212 16882 37268 16884
rect 37212 16830 37214 16882
rect 37214 16830 37266 16882
rect 37266 16830 37268 16882
rect 37212 16828 37268 16830
rect 37996 18396 38052 18452
rect 38108 18226 38164 18228
rect 38108 18174 38110 18226
rect 38110 18174 38162 18226
rect 38162 18174 38164 18226
rect 38108 18172 38164 18174
rect 39676 18844 39732 18900
rect 38892 18450 38948 18452
rect 38892 18398 38894 18450
rect 38894 18398 38946 18450
rect 38946 18398 38948 18450
rect 38892 18396 38948 18398
rect 38556 17724 38612 17780
rect 39676 17500 39732 17556
rect 37996 16994 38052 16996
rect 37996 16942 37998 16994
rect 37998 16942 38050 16994
rect 38050 16942 38052 16994
rect 37996 16940 38052 16942
rect 38892 16268 38948 16324
rect 37436 16156 37492 16212
rect 38332 16210 38388 16212
rect 38332 16158 38334 16210
rect 38334 16158 38386 16210
rect 38386 16158 38388 16210
rect 38332 16156 38388 16158
rect 37324 16098 37380 16100
rect 37324 16046 37326 16098
rect 37326 16046 37378 16098
rect 37378 16046 37380 16098
rect 37324 16044 37380 16046
rect 40012 17276 40068 17332
rect 39788 16828 39844 16884
rect 37324 15820 37380 15876
rect 38892 15538 38948 15540
rect 38892 15486 38894 15538
rect 38894 15486 38946 15538
rect 38946 15486 38948 15538
rect 38892 15484 38948 15486
rect 39564 15484 39620 15540
rect 38108 14812 38164 14868
rect 38892 15036 38948 15092
rect 40124 16492 40180 16548
rect 35980 9772 36036 9828
rect 38892 12962 38948 12964
rect 38892 12910 38894 12962
rect 38894 12910 38946 12962
rect 38946 12910 38948 12962
rect 38892 12908 38948 12910
rect 40012 12850 40068 12852
rect 40012 12798 40014 12850
rect 40014 12798 40066 12850
rect 40066 12798 40068 12850
rect 40012 12796 40068 12798
rect 36428 12684 36484 12740
rect 37100 12738 37156 12740
rect 37100 12686 37102 12738
rect 37102 12686 37154 12738
rect 37154 12686 37156 12738
rect 37100 12684 37156 12686
rect 40124 12124 40180 12180
rect 35868 9042 35924 9044
rect 35868 8990 35870 9042
rect 35870 8990 35922 9042
rect 35922 8990 35924 9042
rect 35868 8988 35924 8990
rect 36428 9042 36484 9044
rect 36428 8990 36430 9042
rect 36430 8990 36482 9042
rect 36482 8990 36484 9042
rect 36428 8988 36484 8990
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 28812 5906 28868 5908
rect 28812 5854 28814 5906
rect 28814 5854 28866 5906
rect 28866 5854 28868 5906
rect 28812 5852 28868 5854
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 32508 5852 32564 5908
rect 38444 5964 38500 6020
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 26124 5346 26180 5348
rect 26124 5294 26126 5346
rect 26126 5294 26178 5346
rect 26178 5294 26180 5346
rect 26124 5292 26180 5294
rect 25788 5234 25844 5236
rect 25788 5182 25790 5234
rect 25790 5182 25842 5234
rect 25842 5182 25844 5234
rect 25788 5180 25844 5182
rect 26348 5180 26404 5236
rect 26236 5122 26292 5124
rect 26236 5070 26238 5122
rect 26238 5070 26290 5122
rect 26290 5070 26292 5122
rect 26236 5068 26292 5070
rect 40124 8092 40180 8148
rect 40012 7420 40068 7476
rect 39676 6748 39732 6804
rect 40124 6076 40180 6132
rect 39788 6018 39844 6020
rect 39788 5966 39790 6018
rect 39790 5966 39842 6018
rect 39842 5966 39844 6018
rect 39788 5964 39844 5966
rect 39564 5906 39620 5908
rect 39564 5854 39566 5906
rect 39566 5854 39618 5906
rect 39618 5854 39620 5906
rect 39564 5852 39620 5854
rect 40124 5906 40180 5908
rect 40124 5854 40126 5906
rect 40126 5854 40178 5906
rect 40178 5854 40180 5906
rect 40124 5852 40180 5854
rect 40124 5404 40180 5460
rect 40124 4732 40180 4788
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 21196 3666 21252 3668
rect 21196 3614 21198 3666
rect 21198 3614 21250 3666
rect 21250 3614 21252 3666
rect 21196 3612 21252 3614
rect 20748 3554 20804 3556
rect 20748 3502 20750 3554
rect 20750 3502 20802 3554
rect 20802 3502 20804 3554
rect 20748 3500 20804 3502
rect 20188 3442 20244 3444
rect 20188 3390 20190 3442
rect 20190 3390 20242 3442
rect 20242 3390 20244 3442
rect 20188 3388 20244 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 40124 4060 40180 4116
rect 40124 3330 40180 3332
rect 40124 3278 40126 3330
rect 40126 3278 40178 3330
rect 40178 3278 40180 3330
rect 40124 3276 40180 3278
rect 39676 2716 39732 2772
rect 39228 2044 39284 2100
<< metal3 >>
rect 41101 43092 41901 43120
rect 38770 43036 38780 43092
rect 38836 43036 41901 43092
rect 41101 43008 41901 43036
rect 41101 42420 41901 42448
rect 40114 42364 40124 42420
rect 40180 42364 41901 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 41101 42336 41901 42364
rect 41101 41748 41901 41776
rect 39218 41692 39228 41748
rect 39284 41692 41901 41748
rect 41101 41664 41901 41692
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 41101 41076 41901 41104
rect 39666 41020 39676 41076
rect 39732 41020 41901 41076
rect 41101 40992 41901 41020
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 0 40404 800 40432
rect 41101 40404 41901 40432
rect 0 40348 1708 40404
rect 1764 40348 1774 40404
rect 25890 40348 25900 40404
rect 25956 40348 26796 40404
rect 26852 40348 29148 40404
rect 29204 40348 29596 40404
rect 29652 40348 29662 40404
rect 40338 40348 40348 40404
rect 40404 40348 41901 40404
rect 0 40320 800 40348
rect 41101 40320 41901 40348
rect 26562 40236 26572 40292
rect 26628 40236 27244 40292
rect 27300 40236 27310 40292
rect 30370 40236 30380 40292
rect 30436 40236 31948 40292
rect 32004 40236 32014 40292
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 0 39732 800 39760
rect 41101 39732 41901 39760
rect 0 39676 4284 39732
rect 4340 39676 4350 39732
rect 40114 39676 40124 39732
rect 40180 39676 41901 39732
rect 0 39648 800 39676
rect 41101 39648 41901 39676
rect 24210 39452 24220 39508
rect 24276 39452 25340 39508
rect 25396 39452 25406 39508
rect 25554 39452 25564 39508
rect 25620 39452 27356 39508
rect 27412 39452 32060 39508
rect 32116 39452 32126 39508
rect 23538 39340 23548 39396
rect 23604 39340 26796 39396
rect 26852 39340 26862 39396
rect 29810 39340 29820 39396
rect 29876 39340 31276 39396
rect 31332 39340 31342 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 41101 39060 41901 39088
rect 40338 39004 40348 39060
rect 40404 39004 41901 39060
rect 41101 38976 41901 39004
rect 30930 38892 30940 38948
rect 30996 38892 32060 38948
rect 32116 38892 32732 38948
rect 32788 38892 32798 38948
rect 23202 38780 23212 38836
rect 23268 38780 25564 38836
rect 25620 38780 25630 38836
rect 28242 38780 28252 38836
rect 28308 38780 30156 38836
rect 30212 38780 30222 38836
rect 27906 38668 27916 38724
rect 27972 38668 29932 38724
rect 29988 38668 29998 38724
rect 31714 38668 31724 38724
rect 31780 38668 33180 38724
rect 33236 38668 33246 38724
rect 29932 38500 29988 38668
rect 30258 38556 30268 38612
rect 30324 38556 31612 38612
rect 31668 38556 31678 38612
rect 29932 38444 31500 38500
rect 31556 38444 31566 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 41101 38388 41901 38416
rect 40114 38332 40124 38388
rect 40180 38332 41901 38388
rect 41101 38304 41901 38332
rect 30146 38108 30156 38164
rect 30212 38108 31052 38164
rect 31108 38108 31118 38164
rect 27906 37996 27916 38052
rect 27972 37996 30828 38052
rect 30884 37996 30894 38052
rect 21410 37884 21420 37940
rect 21476 37884 23212 37940
rect 23268 37884 23278 37940
rect 25106 37884 25116 37940
rect 25172 37884 26572 37940
rect 26628 37884 26638 37940
rect 27346 37884 27356 37940
rect 27412 37884 28588 37940
rect 28644 37884 29540 37940
rect 29698 37884 29708 37940
rect 29764 37884 30492 37940
rect 30548 37884 30558 37940
rect 29484 37828 29540 37884
rect 8418 37772 8428 37828
rect 8484 37772 9660 37828
rect 9716 37772 12460 37828
rect 12516 37772 13356 37828
rect 13412 37772 13422 37828
rect 15810 37772 15820 37828
rect 15876 37772 16716 37828
rect 16772 37772 17612 37828
rect 17668 37772 17678 37828
rect 28130 37772 28140 37828
rect 28196 37772 29148 37828
rect 29204 37772 29214 37828
rect 29484 37772 30268 37828
rect 30324 37772 30334 37828
rect 30594 37772 30604 37828
rect 30660 37772 32172 37828
rect 32228 37772 32238 37828
rect 32498 37772 32508 37828
rect 32564 37772 33292 37828
rect 33348 37772 33358 37828
rect 41101 37716 41901 37744
rect 40114 37660 40124 37716
rect 40180 37660 41901 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 41101 37632 41901 37660
rect 13682 37436 13692 37492
rect 13748 37436 15260 37492
rect 15316 37436 15326 37492
rect 13234 37324 13244 37380
rect 13300 37324 14140 37380
rect 14196 37324 15316 37380
rect 30370 37324 30380 37380
rect 30436 37324 31500 37380
rect 31556 37324 32060 37380
rect 32116 37324 32126 37380
rect 15260 37268 15316 37324
rect 15260 37212 15484 37268
rect 15540 37212 15550 37268
rect 16370 37212 16380 37268
rect 16436 37212 17388 37268
rect 17444 37212 17454 37268
rect 29138 37212 29148 37268
rect 29204 37212 30268 37268
rect 30324 37212 31052 37268
rect 31108 37212 31118 37268
rect 31714 37212 31724 37268
rect 31780 37212 32508 37268
rect 32564 37212 32574 37268
rect 14802 37100 14812 37156
rect 14868 37100 16156 37156
rect 16212 37100 17836 37156
rect 17892 37100 17902 37156
rect 25666 37100 25676 37156
rect 25732 37100 27916 37156
rect 27972 37100 27982 37156
rect 0 37044 800 37072
rect 41101 37044 41901 37072
rect 0 36988 1708 37044
rect 1764 36988 1774 37044
rect 8194 36988 8204 37044
rect 8260 36988 9548 37044
rect 9604 36988 9614 37044
rect 13458 36988 13468 37044
rect 13524 36988 15596 37044
rect 15652 36988 15662 37044
rect 16482 36988 16492 37044
rect 16548 36988 17276 37044
rect 17332 36988 17342 37044
rect 19842 36988 19852 37044
rect 19908 36988 22540 37044
rect 22596 36988 23436 37044
rect 23492 36988 23502 37044
rect 31378 36988 31388 37044
rect 31444 36988 32396 37044
rect 32452 36988 32844 37044
rect 32900 36988 32910 37044
rect 40114 36988 40124 37044
rect 40180 36988 41901 37044
rect 0 36960 800 36988
rect 14812 36932 14868 36988
rect 41101 36960 41901 36988
rect 14802 36876 14812 36932
rect 14868 36876 14878 36932
rect 26114 36876 26124 36932
rect 26180 36876 26460 36932
rect 26516 36876 26526 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 9874 36540 9884 36596
rect 9940 36540 12124 36596
rect 12180 36540 12190 36596
rect 12674 36540 12684 36596
rect 12740 36540 13804 36596
rect 13860 36540 13870 36596
rect 26450 36540 26460 36596
rect 26516 36540 29148 36596
rect 29204 36540 29708 36596
rect 29764 36540 29774 36596
rect 12002 36428 12012 36484
rect 12068 36428 14028 36484
rect 14084 36428 15484 36484
rect 15540 36428 15550 36484
rect 16034 36428 16044 36484
rect 16100 36428 17836 36484
rect 17892 36428 17902 36484
rect 20962 36428 20972 36484
rect 21028 36428 21756 36484
rect 21812 36428 21822 36484
rect 0 36372 800 36400
rect 0 36316 1708 36372
rect 1764 36316 1774 36372
rect 12674 36316 12684 36372
rect 12740 36316 13580 36372
rect 13636 36316 21868 36372
rect 21924 36316 23324 36372
rect 23380 36316 24668 36372
rect 24724 36316 24734 36372
rect 0 36288 800 36316
rect 9762 36204 9772 36260
rect 9828 36204 12460 36260
rect 12516 36204 12526 36260
rect 13906 36204 13916 36260
rect 13972 36204 13982 36260
rect 27234 36204 27244 36260
rect 27300 36204 28476 36260
rect 28532 36204 30380 36260
rect 30436 36204 31276 36260
rect 31332 36204 31342 36260
rect 13916 36148 13972 36204
rect 13916 36092 15148 36148
rect 15204 36092 15596 36148
rect 15652 36092 15662 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 10434 35756 10444 35812
rect 10500 35756 11676 35812
rect 11732 35756 15708 35812
rect 15764 35756 18956 35812
rect 19012 35756 19022 35812
rect 31490 35756 31500 35812
rect 31556 35756 31836 35812
rect 31892 35756 32284 35812
rect 32340 35756 32350 35812
rect 11218 35644 11228 35700
rect 11284 35644 12236 35700
rect 12292 35644 12302 35700
rect 16482 35644 16492 35700
rect 16548 35644 16828 35700
rect 16884 35644 16894 35700
rect 19394 35644 19404 35700
rect 19460 35644 20412 35700
rect 20468 35644 20478 35700
rect 31266 35644 31276 35700
rect 31332 35644 32508 35700
rect 32564 35644 33068 35700
rect 33124 35644 33134 35700
rect 6962 35532 6972 35588
rect 7028 35532 8204 35588
rect 8260 35532 8876 35588
rect 8932 35532 8942 35588
rect 22978 35532 22988 35588
rect 23044 35532 23548 35588
rect 23604 35532 23614 35588
rect 24770 35532 24780 35588
rect 24836 35532 26796 35588
rect 26852 35532 26908 35588
rect 26964 35532 26974 35588
rect 14018 35420 14028 35476
rect 14084 35420 16156 35476
rect 16212 35420 16222 35476
rect 31154 35420 31164 35476
rect 31220 35420 32172 35476
rect 32228 35420 32238 35476
rect 10770 35308 10780 35364
rect 10836 35308 11676 35364
rect 11732 35308 13468 35364
rect 13524 35308 13534 35364
rect 17462 35308 17500 35364
rect 17556 35308 18060 35364
rect 18116 35308 25788 35364
rect 25844 35308 25854 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 26674 35196 26684 35252
rect 26740 35196 27692 35252
rect 27748 35196 27758 35252
rect 31042 35084 31052 35140
rect 31108 35084 31164 35140
rect 31220 35084 31230 35140
rect 15698 34748 15708 34804
rect 15764 34748 16268 34804
rect 16324 34748 19404 34804
rect 19460 34748 19470 34804
rect 30482 34748 30492 34804
rect 30548 34748 31164 34804
rect 31220 34748 31230 34804
rect 10210 34636 10220 34692
rect 10276 34636 11564 34692
rect 11620 34636 13580 34692
rect 13636 34636 15148 34692
rect 15204 34636 15214 34692
rect 17612 34636 23436 34692
rect 23492 34636 23502 34692
rect 28578 34636 28588 34692
rect 28644 34636 29932 34692
rect 29988 34636 31276 34692
rect 31332 34636 31342 34692
rect 17612 34580 17668 34636
rect 12002 34524 12012 34580
rect 12068 34524 14924 34580
rect 14980 34524 14990 34580
rect 15092 34524 16380 34580
rect 16436 34524 17612 34580
rect 17668 34524 17678 34580
rect 30118 34524 30156 34580
rect 30212 34524 30222 34580
rect 15092 34468 15148 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 10892 34412 15148 34468
rect 15250 34412 15260 34468
rect 15316 34412 15326 34468
rect 10892 34244 10948 34412
rect 15260 34356 15316 34412
rect 15260 34300 16604 34356
rect 16660 34300 20188 34356
rect 20244 34300 20254 34356
rect 30482 34300 30492 34356
rect 30548 34300 31052 34356
rect 31108 34300 31118 34356
rect 31266 34300 31276 34356
rect 31332 34300 32396 34356
rect 32452 34300 32462 34356
rect 10882 34188 10892 34244
rect 10948 34188 10958 34244
rect 14914 34188 14924 34244
rect 14980 34188 16044 34244
rect 16100 34188 16110 34244
rect 16482 34188 16492 34244
rect 16548 34188 19516 34244
rect 19572 34188 19852 34244
rect 19908 34188 20524 34244
rect 20580 34188 20590 34244
rect 9650 34076 9660 34132
rect 9716 34076 9726 34132
rect 10994 34076 11004 34132
rect 11060 34076 12124 34132
rect 12180 34076 12190 34132
rect 15474 34076 15484 34132
rect 15540 34076 16604 34132
rect 16660 34076 16670 34132
rect 19730 34076 19740 34132
rect 19796 34076 20300 34132
rect 20356 34076 20366 34132
rect 24098 34076 24108 34132
rect 24164 34076 25452 34132
rect 25508 34076 26236 34132
rect 26292 34076 26302 34132
rect 29250 34076 29260 34132
rect 29316 34076 30156 34132
rect 30212 34076 30222 34132
rect 30482 34076 30492 34132
rect 30548 34076 30940 34132
rect 30996 34076 32284 34132
rect 32340 34076 32350 34132
rect 9660 34020 9716 34076
rect 16604 34020 16660 34076
rect 9202 33964 9212 34020
rect 9268 33964 10892 34020
rect 10948 33964 10958 34020
rect 13794 33964 13804 34020
rect 13860 33964 16380 34020
rect 16436 33964 16446 34020
rect 16604 33964 21532 34020
rect 21588 33964 21598 34020
rect 10658 33852 10668 33908
rect 10724 33852 11340 33908
rect 11396 33852 11406 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 10658 33628 10668 33684
rect 10724 33628 11564 33684
rect 11620 33628 11630 33684
rect 16146 33516 16156 33572
rect 16212 33516 18620 33572
rect 18676 33516 19292 33572
rect 19348 33516 19358 33572
rect 30370 33516 30380 33572
rect 30436 33516 32172 33572
rect 32228 33516 32238 33572
rect 5618 33404 5628 33460
rect 5684 33404 8764 33460
rect 8820 33404 9660 33460
rect 9716 33404 9726 33460
rect 14802 33404 14812 33460
rect 14868 33404 15260 33460
rect 15316 33404 15326 33460
rect 23090 33404 23100 33460
rect 23156 33404 25116 33460
rect 25172 33404 28476 33460
rect 28532 33404 28542 33460
rect 30146 33404 30156 33460
rect 30212 33404 32284 33460
rect 32340 33404 32350 33460
rect 16034 33292 16044 33348
rect 16100 33292 17164 33348
rect 17220 33292 17230 33348
rect 29698 33292 29708 33348
rect 29764 33292 30380 33348
rect 30436 33292 33516 33348
rect 33572 33292 34412 33348
rect 34468 33292 34478 33348
rect 7522 33180 7532 33236
rect 7588 33180 8540 33236
rect 8596 33180 11452 33236
rect 11508 33180 12236 33236
rect 12292 33180 12302 33236
rect 17042 33180 17052 33236
rect 17108 33180 18396 33236
rect 18452 33180 19516 33236
rect 19572 33180 19582 33236
rect 27906 33180 27916 33236
rect 27972 33180 30268 33236
rect 30324 33180 30334 33236
rect 31602 33180 31612 33236
rect 31668 33180 34972 33236
rect 35028 33180 35038 33236
rect 35196 33180 35868 33236
rect 35924 33180 35934 33236
rect 35196 33124 35252 33180
rect 29474 33068 29484 33124
rect 29540 33068 31276 33124
rect 31332 33068 31342 33124
rect 31836 33068 35252 33124
rect 35746 33068 35756 33124
rect 35812 33068 37772 33124
rect 37828 33068 37838 33124
rect 8754 32956 8764 33012
rect 8820 32956 10892 33012
rect 10948 32956 11676 33012
rect 11732 32956 15932 33012
rect 15988 32956 15998 33012
rect 28914 32956 28924 33012
rect 28980 32956 30156 33012
rect 30212 32956 31164 33012
rect 31220 32956 31230 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 31836 32900 31892 33068
rect 31826 32844 31836 32900
rect 31892 32844 31902 32900
rect 18946 32732 18956 32788
rect 19012 32732 19740 32788
rect 19796 32732 19806 32788
rect 20626 32732 20636 32788
rect 20692 32732 23212 32788
rect 23268 32732 23278 32788
rect 26002 32732 26012 32788
rect 26068 32732 27356 32788
rect 27412 32732 27422 32788
rect 28130 32732 28140 32788
rect 28196 32732 32172 32788
rect 32228 32732 32238 32788
rect 22978 32620 22988 32676
rect 23044 32620 31612 32676
rect 31668 32620 31678 32676
rect 7634 32508 7644 32564
rect 7700 32508 8204 32564
rect 8260 32508 8270 32564
rect 15810 32508 15820 32564
rect 15876 32508 17388 32564
rect 17444 32508 17454 32564
rect 18386 32508 18396 32564
rect 18452 32508 18844 32564
rect 18900 32508 19404 32564
rect 19460 32508 20636 32564
rect 20692 32508 20702 32564
rect 25778 32508 25788 32564
rect 25844 32508 29036 32564
rect 29092 32508 29102 32564
rect 29250 32508 29260 32564
rect 29316 32508 31500 32564
rect 31556 32508 31566 32564
rect 33180 32508 36652 32564
rect 36708 32508 37100 32564
rect 37156 32508 37166 32564
rect 33180 32452 33236 32508
rect 8082 32396 8092 32452
rect 8148 32396 8652 32452
rect 8708 32396 8718 32452
rect 24658 32396 24668 32452
rect 24724 32396 25564 32452
rect 25620 32396 25630 32452
rect 26002 32396 26012 32452
rect 26068 32396 33236 32452
rect 33394 32396 33404 32452
rect 33460 32396 33964 32452
rect 34020 32396 35644 32452
rect 35700 32396 35710 32452
rect 17714 32284 17724 32340
rect 17780 32284 19068 32340
rect 19124 32284 20300 32340
rect 20356 32284 20366 32340
rect 30034 32284 30044 32340
rect 30100 32284 33628 32340
rect 33684 32284 34188 32340
rect 34244 32284 34254 32340
rect 30818 32172 30828 32228
rect 30884 32172 31388 32228
rect 31444 32172 31454 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 10098 31948 10108 32004
rect 10164 31948 11676 32004
rect 11732 31948 17164 32004
rect 17220 31948 17230 32004
rect 36418 31948 36428 32004
rect 36484 31948 36876 32004
rect 36932 31948 36942 32004
rect 15138 31836 15148 31892
rect 15204 31836 15820 31892
rect 15876 31836 15886 31892
rect 16930 31836 16940 31892
rect 16996 31836 18956 31892
rect 19012 31836 19022 31892
rect 19842 31836 19852 31892
rect 19908 31836 20748 31892
rect 20804 31836 20814 31892
rect 23538 31836 23548 31892
rect 23604 31836 27020 31892
rect 27076 31836 27580 31892
rect 27636 31836 27646 31892
rect 27794 31836 27804 31892
rect 27860 31836 29596 31892
rect 29652 31836 29662 31892
rect 34626 31836 34636 31892
rect 34692 31836 36764 31892
rect 36820 31836 36830 31892
rect 36978 31836 36988 31892
rect 37044 31836 37884 31892
rect 37940 31836 37950 31892
rect 27804 31780 27860 31836
rect 16594 31724 16604 31780
rect 16660 31724 18172 31780
rect 18228 31724 18508 31780
rect 18564 31724 18574 31780
rect 20066 31724 20076 31780
rect 20132 31724 21420 31780
rect 21476 31724 21486 31780
rect 22418 31724 22428 31780
rect 22484 31724 23324 31780
rect 23380 31724 24108 31780
rect 24164 31724 26236 31780
rect 26292 31724 26302 31780
rect 26562 31724 26572 31780
rect 26628 31724 27860 31780
rect 31826 31724 31836 31780
rect 31892 31724 35756 31780
rect 35812 31724 35822 31780
rect 35970 31724 35980 31780
rect 36036 31724 37100 31780
rect 37156 31724 37166 31780
rect 11442 31612 11452 31668
rect 11508 31612 12684 31668
rect 12740 31612 12750 31668
rect 15092 31612 24668 31668
rect 24724 31612 24734 31668
rect 25330 31612 25340 31668
rect 25396 31612 30156 31668
rect 30212 31612 30222 31668
rect 36530 31612 36540 31668
rect 36596 31612 37548 31668
rect 37604 31612 37614 31668
rect 15092 31556 15148 31612
rect 9202 31500 9212 31556
rect 9268 31500 15148 31556
rect 21522 31500 21532 31556
rect 21588 31500 23548 31556
rect 23604 31500 23614 31556
rect 23874 31500 23884 31556
rect 23940 31500 25004 31556
rect 25060 31500 25070 31556
rect 26786 31500 26796 31556
rect 26852 31500 28028 31556
rect 28084 31500 29820 31556
rect 29876 31500 29886 31556
rect 35298 31500 35308 31556
rect 35364 31500 36316 31556
rect 36372 31500 37212 31556
rect 37268 31500 37278 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 26226 31276 26236 31332
rect 26292 31276 26908 31332
rect 34178 31276 34188 31332
rect 34244 31276 36316 31332
rect 36372 31276 36382 31332
rect 26852 31220 26908 31276
rect 8306 31164 8316 31220
rect 8372 31164 22204 31220
rect 22260 31164 22988 31220
rect 23044 31164 23054 31220
rect 26852 31164 35868 31220
rect 35924 31164 35934 31220
rect 26226 31052 26236 31108
rect 26292 31052 26302 31108
rect 30146 31052 30156 31108
rect 30212 31052 35084 31108
rect 35140 31052 35150 31108
rect 26236 30996 26292 31052
rect 18946 30940 18956 30996
rect 19012 30940 24332 30996
rect 24388 30940 25676 30996
rect 25732 30940 26292 30996
rect 16370 30828 16380 30884
rect 16436 30828 17500 30884
rect 17556 30828 17566 30884
rect 23762 30828 23772 30884
rect 23828 30828 30716 30884
rect 30772 30828 30782 30884
rect 35634 30828 35644 30884
rect 35700 30828 37660 30884
rect 37716 30828 37726 30884
rect 18274 30716 18284 30772
rect 18340 30716 19068 30772
rect 19124 30716 19134 30772
rect 26002 30716 26012 30772
rect 26068 30716 26572 30772
rect 26628 30716 26638 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 24658 30492 24668 30548
rect 24724 30492 26572 30548
rect 26628 30492 26638 30548
rect 26852 30492 28364 30548
rect 28420 30492 29484 30548
rect 29540 30492 31164 30548
rect 31220 30492 31230 30548
rect 26852 30324 26908 30492
rect 5954 30268 5964 30324
rect 6020 30268 8204 30324
rect 8260 30268 8270 30324
rect 22194 30268 22204 30324
rect 22260 30268 22988 30324
rect 23044 30268 24108 30324
rect 24164 30268 24174 30324
rect 24546 30268 24556 30324
rect 24612 30268 26908 30324
rect 28476 30268 30604 30324
rect 30660 30268 30670 30324
rect 30818 30268 30828 30324
rect 30884 30268 32060 30324
rect 32116 30268 32126 30324
rect 34626 30268 34636 30324
rect 34692 30268 35868 30324
rect 35924 30268 35934 30324
rect 38612 30268 40124 30324
rect 40180 30268 40190 30324
rect 8866 30156 8876 30212
rect 8932 30156 9884 30212
rect 9940 30156 9950 30212
rect 16706 30156 16716 30212
rect 16772 30156 17948 30212
rect 18004 30156 18732 30212
rect 18788 30156 18798 30212
rect 25778 30156 25788 30212
rect 25844 30156 26460 30212
rect 26516 30156 26526 30212
rect 26786 30156 26796 30212
rect 26852 30156 27132 30212
rect 27188 30156 27198 30212
rect 20850 30044 20860 30100
rect 20916 30044 21868 30100
rect 21924 30044 21934 30100
rect 26460 29988 26516 30156
rect 28476 30100 28532 30268
rect 38612 30212 38668 30268
rect 32162 30156 32172 30212
rect 32228 30156 32732 30212
rect 32788 30156 32798 30212
rect 32946 30156 32956 30212
rect 33012 30156 33964 30212
rect 34020 30156 34030 30212
rect 36194 30156 36204 30212
rect 36260 30156 37324 30212
rect 37380 30156 38668 30212
rect 26898 30044 26908 30100
rect 26964 30044 28252 30100
rect 28308 30044 28532 30100
rect 29586 30044 29596 30100
rect 29652 30044 30044 30100
rect 30100 30044 30380 30100
rect 30436 30044 34524 30100
rect 34580 30044 34590 30100
rect 26908 29988 26964 30044
rect 7522 29932 7532 29988
rect 7588 29932 8316 29988
rect 8372 29932 10108 29988
rect 10164 29932 10174 29988
rect 18498 29932 18508 29988
rect 18564 29932 19404 29988
rect 19460 29932 19470 29988
rect 21522 29932 21532 29988
rect 21588 29932 22764 29988
rect 22820 29932 22830 29988
rect 26460 29932 26964 29988
rect 27122 29932 27132 29988
rect 27188 29932 29148 29988
rect 29204 29932 29214 29988
rect 30258 29932 30268 29988
rect 30324 29932 35980 29988
rect 36036 29932 36876 29988
rect 36932 29932 36942 29988
rect 37874 29932 37884 29988
rect 37940 29932 38444 29988
rect 38500 29932 38510 29988
rect 16706 29820 16716 29876
rect 16772 29820 19180 29876
rect 19236 29820 19246 29876
rect 29250 29820 29260 29876
rect 29316 29820 30380 29876
rect 30436 29820 31836 29876
rect 31892 29820 31902 29876
rect 32834 29820 32844 29876
rect 32900 29820 34076 29876
rect 34132 29820 34142 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 30594 29708 30604 29764
rect 30660 29708 31948 29764
rect 32004 29708 33292 29764
rect 33348 29708 33358 29764
rect 16146 29596 16156 29652
rect 16212 29596 16716 29652
rect 16772 29596 18396 29652
rect 18452 29596 18462 29652
rect 26852 29596 28308 29652
rect 28466 29596 28476 29652
rect 28532 29596 30492 29652
rect 30548 29596 32396 29652
rect 32452 29596 32462 29652
rect 26852 29540 26908 29596
rect 28252 29540 28308 29596
rect 16930 29484 16940 29540
rect 16996 29484 17500 29540
rect 17556 29484 17566 29540
rect 23314 29484 23324 29540
rect 23380 29484 25116 29540
rect 25172 29484 26908 29540
rect 27010 29484 27020 29540
rect 27076 29484 27086 29540
rect 28252 29484 37884 29540
rect 37940 29484 37950 29540
rect 27020 29428 27076 29484
rect 8642 29372 8652 29428
rect 8708 29372 9436 29428
rect 9492 29372 9772 29428
rect 9828 29372 11116 29428
rect 11172 29372 11182 29428
rect 12226 29372 12236 29428
rect 12292 29372 13580 29428
rect 13636 29372 13646 29428
rect 15698 29372 15708 29428
rect 15764 29372 17388 29428
rect 17444 29372 17454 29428
rect 20402 29372 20412 29428
rect 20468 29372 21420 29428
rect 21476 29372 21486 29428
rect 26562 29372 26572 29428
rect 26628 29372 27076 29428
rect 30818 29372 30828 29428
rect 30884 29372 31500 29428
rect 31556 29372 33628 29428
rect 33684 29372 35644 29428
rect 35700 29372 35710 29428
rect 35858 29372 35868 29428
rect 35924 29372 38220 29428
rect 38276 29372 38286 29428
rect 7074 29260 7084 29316
rect 7140 29260 9996 29316
rect 10052 29260 10062 29316
rect 12898 29260 12908 29316
rect 12964 29260 13916 29316
rect 13972 29260 13982 29316
rect 21074 29260 21084 29316
rect 21140 29260 21868 29316
rect 21924 29260 21934 29316
rect 38546 29260 38556 29316
rect 38612 29260 40124 29316
rect 40180 29260 40190 29316
rect 10322 29148 10332 29204
rect 10388 29148 10780 29204
rect 10836 29148 10846 29204
rect 11666 29148 11676 29204
rect 11732 29148 16156 29204
rect 16212 29148 16222 29204
rect 17490 29148 17500 29204
rect 17556 29148 19852 29204
rect 19908 29148 19918 29204
rect 33842 29148 33852 29204
rect 33908 29148 35532 29204
rect 35588 29148 35598 29204
rect 13794 29036 13804 29092
rect 13860 29036 18060 29092
rect 18116 29036 19628 29092
rect 19684 29036 19694 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 10098 28924 10108 28980
rect 10164 28924 10444 28980
rect 10500 28924 12124 28980
rect 12180 28924 12190 28980
rect 11106 28812 11116 28868
rect 11172 28812 12460 28868
rect 12516 28812 12526 28868
rect 17490 28812 17500 28868
rect 17556 28812 18844 28868
rect 18900 28812 18910 28868
rect 9202 28700 9212 28756
rect 9268 28700 9884 28756
rect 9940 28700 12572 28756
rect 12628 28700 12638 28756
rect 24658 28700 24668 28756
rect 24724 28700 25228 28756
rect 25284 28700 28476 28756
rect 28532 28700 30268 28756
rect 30324 28700 30940 28756
rect 30996 28700 31006 28756
rect 4722 28588 4732 28644
rect 4788 28588 6300 28644
rect 6356 28588 6366 28644
rect 11554 28588 11564 28644
rect 11620 28588 12348 28644
rect 12404 28588 12796 28644
rect 12852 28588 12862 28644
rect 16146 28588 16156 28644
rect 16212 28588 18172 28644
rect 18228 28588 18238 28644
rect 31266 28588 31276 28644
rect 31332 28588 32172 28644
rect 32228 28588 32238 28644
rect 12002 28476 12012 28532
rect 12068 28476 13468 28532
rect 13524 28476 13534 28532
rect 26898 28476 26908 28532
rect 26964 28476 27916 28532
rect 27972 28476 27982 28532
rect 12898 28364 12908 28420
rect 12964 28364 13580 28420
rect 13636 28364 13646 28420
rect 23650 28364 23660 28420
rect 23716 28364 24780 28420
rect 24836 28364 24846 28420
rect 34402 28364 34412 28420
rect 34468 28364 35532 28420
rect 35588 28364 35598 28420
rect 24098 28252 24108 28308
rect 24164 28252 25452 28308
rect 25508 28252 25788 28308
rect 25844 28252 25854 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 14130 28028 14140 28084
rect 14196 28028 17500 28084
rect 17556 28028 17566 28084
rect 32284 28028 33068 28084
rect 33124 28028 33134 28084
rect 32284 27972 32340 28028
rect 27346 27916 27356 27972
rect 27412 27916 32284 27972
rect 32340 27916 32350 27972
rect 9538 27804 9548 27860
rect 9604 27804 9614 27860
rect 15922 27804 15932 27860
rect 15988 27804 16380 27860
rect 16436 27804 23324 27860
rect 23380 27804 27244 27860
rect 27300 27804 27310 27860
rect 27906 27804 27916 27860
rect 27972 27804 29036 27860
rect 29092 27804 29102 27860
rect 32050 27804 32060 27860
rect 32116 27804 33852 27860
rect 33908 27804 33918 27860
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 9548 27412 9604 27804
rect 18722 27692 18732 27748
rect 18788 27692 19404 27748
rect 19460 27692 19470 27748
rect 29810 27580 29820 27636
rect 29876 27580 31948 27636
rect 32004 27580 32014 27636
rect 33292 27580 35420 27636
rect 35476 27580 35486 27636
rect 33292 27524 33348 27580
rect 32050 27468 32060 27524
rect 32116 27468 33348 27524
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 9426 27356 9436 27412
rect 9492 27356 10556 27412
rect 10612 27356 23772 27412
rect 23828 27356 24332 27412
rect 24388 27356 25340 27412
rect 25396 27356 25406 27412
rect 31154 27356 31164 27412
rect 31220 27356 32284 27412
rect 32340 27356 32350 27412
rect 6962 27244 6972 27300
rect 7028 27244 22540 27300
rect 22596 27244 22606 27300
rect 33506 27244 33516 27300
rect 33572 27244 35308 27300
rect 35364 27244 35374 27300
rect 36306 27244 36316 27300
rect 36372 27244 37996 27300
rect 38052 27244 38062 27300
rect 36316 27188 36372 27244
rect 16706 27132 16716 27188
rect 16772 27132 18508 27188
rect 18564 27132 18574 27188
rect 19282 27132 19292 27188
rect 19348 27132 21308 27188
rect 21364 27132 21374 27188
rect 30034 27132 30044 27188
rect 30100 27132 31612 27188
rect 31668 27132 31678 27188
rect 34850 27132 34860 27188
rect 34916 27132 36372 27188
rect 19628 27020 20412 27076
rect 20468 27020 20478 27076
rect 23538 27020 23548 27076
rect 23604 27020 24108 27076
rect 24164 27020 29596 27076
rect 29652 27020 29662 27076
rect 31714 27020 31724 27076
rect 31780 27020 32900 27076
rect 34738 27020 34748 27076
rect 34804 27020 35420 27076
rect 35476 27020 35486 27076
rect 3938 26908 3948 26964
rect 4004 26908 5628 26964
rect 5684 26908 6188 26964
rect 6244 26908 6254 26964
rect 14242 26908 14252 26964
rect 14308 26908 17780 26964
rect 17724 26852 17780 26908
rect 19628 26852 19684 27020
rect 20738 26908 20748 26964
rect 20804 26908 23436 26964
rect 23492 26908 23502 26964
rect 27570 26908 27580 26964
rect 27636 26908 28588 26964
rect 28644 26908 28654 26964
rect 29922 26908 29932 26964
rect 29988 26908 31388 26964
rect 31444 26908 31454 26964
rect 32844 26852 32900 27020
rect 41101 26964 41901 26992
rect 33058 26908 33068 26964
rect 33124 26908 33740 26964
rect 33796 26908 34524 26964
rect 34580 26908 34590 26964
rect 40124 26908 41901 26964
rect 34524 26852 34580 26908
rect 40124 26852 40180 26908
rect 41101 26880 41901 26908
rect 17714 26796 17724 26852
rect 17780 26796 17790 26852
rect 19618 26796 19628 26852
rect 19684 26796 19694 26852
rect 28354 26796 28364 26852
rect 28420 26796 29484 26852
rect 29540 26796 29550 26852
rect 32834 26796 32844 26852
rect 32900 26796 32910 26852
rect 34524 26796 36316 26852
rect 36372 26796 36382 26852
rect 39554 26796 39564 26852
rect 39620 26796 40124 26852
rect 40180 26796 40190 26852
rect 19394 26684 19404 26740
rect 19460 26684 19470 26740
rect 17602 26460 17612 26516
rect 17668 26460 18396 26516
rect 18452 26460 19180 26516
rect 19236 26460 19246 26516
rect 19404 26404 19460 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 24322 26572 24332 26628
rect 24388 26572 39788 26628
rect 39844 26572 39854 26628
rect 32610 26460 32620 26516
rect 32676 26460 33292 26516
rect 33348 26460 33358 26516
rect 19058 26348 19068 26404
rect 19124 26348 19460 26404
rect 41101 26292 41901 26320
rect 27682 26236 27692 26292
rect 27748 26236 30940 26292
rect 30996 26236 31006 26292
rect 32050 26236 32060 26292
rect 32116 26236 33292 26292
rect 33348 26236 33358 26292
rect 40002 26236 40012 26292
rect 40068 26236 41901 26292
rect 41101 26208 41901 26236
rect 26226 26124 26236 26180
rect 26292 26124 26908 26180
rect 26964 26124 27524 26180
rect 28242 26124 28252 26180
rect 28308 26124 35308 26180
rect 35364 26124 35374 26180
rect 27468 26068 27524 26124
rect 27468 26012 28588 26068
rect 28644 26012 28654 26068
rect 31490 26012 31500 26068
rect 31556 26012 32732 26068
rect 32788 26012 32798 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 10770 25564 10780 25620
rect 10836 25564 11452 25620
rect 11508 25564 14140 25620
rect 14196 25564 14206 25620
rect 31126 25564 31164 25620
rect 31220 25564 31230 25620
rect 23874 25452 23884 25508
rect 23940 25452 24780 25508
rect 24836 25452 24846 25508
rect 30258 25452 30268 25508
rect 30324 25452 30828 25508
rect 30884 25452 30894 25508
rect 2034 25340 2044 25396
rect 2100 25340 10220 25396
rect 10276 25340 10892 25396
rect 10948 25340 10958 25396
rect 22754 25340 22764 25396
rect 22820 25340 23212 25396
rect 23268 25340 23772 25396
rect 23828 25340 23838 25396
rect 24210 25340 24220 25396
rect 24276 25340 26908 25396
rect 31602 25340 31612 25396
rect 31668 25340 32172 25396
rect 32228 25340 33852 25396
rect 33908 25340 33918 25396
rect 26852 25284 26908 25340
rect 8642 25228 8652 25284
rect 8708 25228 9212 25284
rect 9268 25228 11004 25284
rect 11060 25228 21532 25284
rect 21588 25228 21598 25284
rect 26852 25228 39788 25284
rect 39844 25228 39854 25284
rect 1698 25116 1708 25172
rect 1764 25116 2940 25172
rect 2996 25116 5068 25172
rect 5124 25116 5134 25172
rect 32946 25116 32956 25172
rect 33012 25116 33292 25172
rect 33348 25116 33358 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 4162 25004 4172 25060
rect 4228 25004 6412 25060
rect 6468 25004 6478 25060
rect 11106 25004 11116 25060
rect 11172 25004 18508 25060
rect 18564 25004 18574 25060
rect 0 24948 800 24976
rect 0 24892 1708 24948
rect 1764 24892 2492 24948
rect 2548 24892 2558 24948
rect 0 24864 800 24892
rect 5282 24780 5292 24836
rect 5348 24780 6412 24836
rect 6468 24780 6478 24836
rect 10322 24780 10332 24836
rect 10388 24780 10892 24836
rect 10948 24780 14028 24836
rect 14084 24780 14094 24836
rect 22306 24780 22316 24836
rect 22372 24780 25564 24836
rect 25620 24780 25630 24836
rect 4610 24668 4620 24724
rect 4676 24668 11564 24724
rect 11620 24668 13356 24724
rect 13412 24668 13422 24724
rect 21186 24668 21196 24724
rect 21252 24668 22092 24724
rect 22148 24668 22158 24724
rect 24994 24668 25004 24724
rect 25060 24668 25788 24724
rect 25844 24668 26684 24724
rect 26740 24668 26750 24724
rect 31378 24668 31388 24724
rect 31444 24668 32956 24724
rect 33012 24668 33022 24724
rect 4162 24556 4172 24612
rect 4228 24556 7532 24612
rect 7588 24556 7598 24612
rect 12338 24556 12348 24612
rect 12404 24556 17612 24612
rect 17668 24556 17678 24612
rect 35746 24556 35756 24612
rect 35812 24556 40124 24612
rect 40180 24556 40190 24612
rect 15092 24332 20636 24388
rect 20692 24332 20702 24388
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 0 24220 1932 24276
rect 1988 24220 1998 24276
rect 0 24192 800 24220
rect 15092 24164 15148 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 2930 24108 2940 24164
rect 2996 24108 15148 24164
rect 17826 24108 17836 24164
rect 17892 24108 17902 24164
rect 20178 24108 20188 24164
rect 20244 24108 20748 24164
rect 20804 24108 20814 24164
rect 17836 23940 17892 24108
rect 18498 23996 18508 24052
rect 18564 23996 18956 24052
rect 19012 23996 23772 24052
rect 23828 23996 25228 24052
rect 25284 23996 25294 24052
rect 34066 23996 34076 24052
rect 34132 23996 36764 24052
rect 36820 23996 40124 24052
rect 40180 23996 40190 24052
rect 6290 23884 6300 23940
rect 6356 23884 7980 23940
rect 8036 23884 8652 23940
rect 8708 23884 8718 23940
rect 11554 23884 11564 23940
rect 11620 23884 12348 23940
rect 12404 23884 12414 23940
rect 16818 23884 16828 23940
rect 16884 23884 17052 23940
rect 17108 23884 17118 23940
rect 17266 23884 17276 23940
rect 17332 23884 18172 23940
rect 18228 23884 18238 23940
rect 19842 23884 19852 23940
rect 19908 23884 21420 23940
rect 21476 23884 21486 23940
rect 23090 23884 23100 23940
rect 23156 23884 24220 23940
rect 24276 23884 24286 23940
rect 36530 23884 36540 23940
rect 36596 23884 37212 23940
rect 37268 23884 37278 23940
rect 14242 23772 14252 23828
rect 14308 23772 18060 23828
rect 18116 23772 18126 23828
rect 20178 23772 20188 23828
rect 20244 23772 22764 23828
rect 22820 23772 22830 23828
rect 4722 23660 4732 23716
rect 4788 23660 6524 23716
rect 6580 23660 6590 23716
rect 16370 23660 16380 23716
rect 16436 23660 16828 23716
rect 16884 23660 16894 23716
rect 18162 23660 18172 23716
rect 18228 23660 20076 23716
rect 20132 23660 20142 23716
rect 21634 23660 21644 23716
rect 21700 23660 22316 23716
rect 22372 23660 22382 23716
rect 16828 23604 16884 23660
rect 8866 23548 8876 23604
rect 8932 23548 9772 23604
rect 9828 23548 9838 23604
rect 16828 23548 19628 23604
rect 19684 23548 19694 23604
rect 32050 23548 32060 23604
rect 32116 23548 33740 23604
rect 33796 23548 33806 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 5282 23436 5292 23492
rect 5348 23436 7420 23492
rect 7476 23436 7486 23492
rect 21298 23436 21308 23492
rect 21364 23436 27804 23492
rect 27860 23436 27870 23492
rect 3266 23324 3276 23380
rect 3332 23324 3836 23380
rect 3892 23324 3902 23380
rect 5170 23324 5180 23380
rect 5236 23324 7196 23380
rect 7252 23324 7644 23380
rect 7700 23324 7710 23380
rect 9874 23324 9884 23380
rect 9940 23324 21868 23380
rect 21924 23324 23100 23380
rect 23156 23324 23166 23380
rect 30482 23324 30492 23380
rect 30548 23324 34188 23380
rect 34244 23324 34254 23380
rect 36642 23324 36652 23380
rect 36708 23324 38332 23380
rect 38388 23324 38398 23380
rect 36652 23268 36708 23324
rect 5058 23212 5068 23268
rect 5124 23212 7420 23268
rect 7476 23212 7486 23268
rect 15446 23212 15484 23268
rect 15540 23212 15550 23268
rect 16370 23212 16380 23268
rect 16436 23212 21308 23268
rect 21364 23212 21374 23268
rect 24434 23212 24444 23268
rect 24500 23212 27468 23268
rect 27524 23212 27534 23268
rect 29138 23212 29148 23268
rect 29204 23212 30044 23268
rect 30100 23212 30110 23268
rect 33730 23212 33740 23268
rect 33796 23212 36708 23268
rect 4386 23100 4396 23156
rect 4452 23100 5628 23156
rect 5684 23100 5694 23156
rect 13010 23100 13020 23156
rect 13076 23100 16268 23156
rect 16324 23100 16334 23156
rect 17938 23100 17948 23156
rect 18004 23100 18508 23156
rect 18564 23100 22092 23156
rect 22148 23100 22158 23156
rect 4274 22988 4284 23044
rect 4340 22988 19068 23044
rect 19124 22988 19516 23044
rect 19572 22988 19582 23044
rect 27794 22988 27804 23044
rect 27860 22988 29932 23044
rect 29988 22988 29998 23044
rect 4498 22876 4508 22932
rect 4564 22876 6636 22932
rect 6692 22876 6702 22932
rect 5618 22764 5628 22820
rect 5684 22764 6412 22820
rect 6468 22764 6478 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 5506 22652 5516 22708
rect 5572 22652 6524 22708
rect 6580 22652 6590 22708
rect 4946 22540 4956 22596
rect 5012 22540 6412 22596
rect 6468 22540 6478 22596
rect 15698 22540 15708 22596
rect 15764 22540 16716 22596
rect 16772 22540 17612 22596
rect 17668 22540 17678 22596
rect 27458 22540 27468 22596
rect 27524 22540 29036 22596
rect 29092 22540 29102 22596
rect 5058 22428 5068 22484
rect 5124 22428 6300 22484
rect 6356 22428 6366 22484
rect 6626 22428 6636 22484
rect 6692 22428 11340 22484
rect 11396 22428 11406 22484
rect 18610 22428 18620 22484
rect 18676 22428 19404 22484
rect 19460 22428 28252 22484
rect 28308 22428 28318 22484
rect 31266 22428 31276 22484
rect 31332 22428 33404 22484
rect 33460 22428 33470 22484
rect 4844 22316 6748 22372
rect 6804 22316 8428 22372
rect 8484 22316 8652 22372
rect 8708 22316 8718 22372
rect 19618 22316 19628 22372
rect 19684 22316 20524 22372
rect 20580 22316 20972 22372
rect 21028 22316 21038 22372
rect 33282 22316 33292 22372
rect 33348 22316 34188 22372
rect 34244 22316 35532 22372
rect 35588 22316 37324 22372
rect 37380 22316 37390 22372
rect 4844 22260 4900 22316
rect 4806 22204 4844 22260
rect 4900 22204 4910 22260
rect 18722 22204 18732 22260
rect 18788 22204 28028 22260
rect 28084 22204 28094 22260
rect 28466 22204 28476 22260
rect 28532 22204 29988 22260
rect 33058 22204 33068 22260
rect 33124 22204 34412 22260
rect 34468 22204 35868 22260
rect 35924 22204 35934 22260
rect 29932 22148 29988 22204
rect 5394 22092 5404 22148
rect 5460 22092 6300 22148
rect 6356 22092 6524 22148
rect 6580 22092 6590 22148
rect 26338 22092 26348 22148
rect 26404 22092 26908 22148
rect 26964 22092 27244 22148
rect 27300 22092 27310 22148
rect 27906 22092 27916 22148
rect 27972 22092 29148 22148
rect 29204 22092 29214 22148
rect 29922 22092 29932 22148
rect 29988 22092 33404 22148
rect 33460 22092 33470 22148
rect 34626 22092 34636 22148
rect 34692 22092 36316 22148
rect 36372 22092 36876 22148
rect 36932 22092 38444 22148
rect 38500 22092 38510 22148
rect 33506 21980 33516 22036
rect 33572 21980 35196 22036
rect 35252 21980 35262 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 6738 21868 6748 21924
rect 6804 21868 7084 21924
rect 7140 21868 7150 21924
rect 14466 21868 14476 21924
rect 14532 21868 16044 21924
rect 16100 21868 16716 21924
rect 16772 21868 16782 21924
rect 22082 21868 22092 21924
rect 22148 21868 23100 21924
rect 23156 21868 23166 21924
rect 1698 21756 1708 21812
rect 1764 21756 3052 21812
rect 3108 21756 3500 21812
rect 3556 21756 3566 21812
rect 5730 21756 5740 21812
rect 5796 21756 7196 21812
rect 7252 21756 7262 21812
rect 11666 21756 11676 21812
rect 11732 21756 15652 21812
rect 17490 21756 17500 21812
rect 17556 21756 18396 21812
rect 18452 21756 18462 21812
rect 26786 21756 26796 21812
rect 26852 21756 29652 21812
rect 36418 21756 36428 21812
rect 36484 21756 37268 21812
rect 5058 21644 5068 21700
rect 5124 21644 5852 21700
rect 5908 21644 5918 21700
rect 6626 21644 6636 21700
rect 6692 21644 7532 21700
rect 7588 21644 7598 21700
rect 12002 21644 12012 21700
rect 12068 21644 13916 21700
rect 13972 21644 15372 21700
rect 15428 21644 15438 21700
rect 15596 21588 15652 21756
rect 29596 21700 29652 21756
rect 37212 21700 37268 21756
rect 17938 21644 17948 21700
rect 18004 21644 19292 21700
rect 19348 21644 19358 21700
rect 29586 21644 29596 21700
rect 29652 21644 29662 21700
rect 31714 21644 31724 21700
rect 31780 21644 34860 21700
rect 34916 21644 35084 21700
rect 35140 21644 35532 21700
rect 35588 21644 35598 21700
rect 36082 21644 36092 21700
rect 36148 21644 36988 21700
rect 37044 21644 37054 21700
rect 37202 21644 37212 21700
rect 37268 21644 38556 21700
rect 38612 21644 38622 21700
rect 3826 21532 3836 21588
rect 3892 21532 4620 21588
rect 4676 21532 4686 21588
rect 15250 21532 15260 21588
rect 15316 21532 16156 21588
rect 16212 21532 18172 21588
rect 18228 21532 19180 21588
rect 19236 21532 19246 21588
rect 27570 21532 27580 21588
rect 27636 21532 28812 21588
rect 28868 21532 28878 21588
rect 32162 21532 32172 21588
rect 32228 21532 32732 21588
rect 32788 21532 33180 21588
rect 33236 21532 33246 21588
rect 33814 21532 33852 21588
rect 33908 21532 33918 21588
rect 35410 21532 35420 21588
rect 35476 21532 38108 21588
rect 38164 21532 40124 21588
rect 40180 21532 40190 21588
rect 6738 21420 6748 21476
rect 6804 21420 7196 21476
rect 7252 21420 7262 21476
rect 15586 21420 15596 21476
rect 15652 21420 21532 21476
rect 21588 21420 21598 21476
rect 23762 21420 23772 21476
rect 23828 21420 24220 21476
rect 24276 21420 25340 21476
rect 25396 21420 25788 21476
rect 25844 21420 26124 21476
rect 26180 21420 26572 21476
rect 26628 21420 26638 21476
rect 33282 21420 33292 21476
rect 33348 21420 34188 21476
rect 34244 21420 34254 21476
rect 13570 21308 13580 21364
rect 13636 21308 15484 21364
rect 15540 21308 16268 21364
rect 16324 21308 16334 21364
rect 17042 21308 17052 21364
rect 17108 21308 18060 21364
rect 18116 21308 19068 21364
rect 19124 21308 19134 21364
rect 29586 21308 29596 21364
rect 29652 21308 37436 21364
rect 37492 21308 37502 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 16818 21084 16828 21140
rect 16884 21084 17388 21140
rect 17444 21084 17454 21140
rect 4946 20972 4956 21028
rect 5012 20972 6188 21028
rect 6244 20972 6254 21028
rect 17714 20972 17724 21028
rect 17780 20972 17948 21028
rect 18004 20972 18014 21028
rect 29810 20972 29820 21028
rect 29876 20972 30828 21028
rect 30884 20972 30894 21028
rect 41101 20916 41901 20944
rect 8978 20860 8988 20916
rect 9044 20860 18844 20916
rect 18900 20860 18910 20916
rect 40002 20860 40012 20916
rect 40068 20860 41901 20916
rect 41101 20832 41901 20860
rect 6066 20748 6076 20804
rect 6132 20748 6636 20804
rect 6692 20748 9548 20804
rect 9604 20748 10108 20804
rect 10164 20748 10174 20804
rect 16370 20748 16380 20804
rect 16436 20748 17276 20804
rect 17332 20748 17836 20804
rect 17892 20748 17902 20804
rect 21746 20748 21756 20804
rect 21812 20748 23884 20804
rect 23940 20748 25788 20804
rect 25844 20748 25854 20804
rect 28130 20748 28140 20804
rect 28196 20748 29484 20804
rect 29540 20748 29550 20804
rect 32498 20748 32508 20804
rect 32564 20748 34188 20804
rect 34244 20748 34254 20804
rect 4722 20636 4732 20692
rect 4788 20636 8540 20692
rect 8596 20636 9212 20692
rect 9268 20636 9278 20692
rect 17154 20636 17164 20692
rect 17220 20636 18172 20692
rect 18228 20636 18238 20692
rect 32610 20636 32620 20692
rect 32676 20636 34748 20692
rect 34804 20636 34814 20692
rect 2370 20524 2380 20580
rect 2436 20524 3612 20580
rect 3668 20524 4172 20580
rect 4228 20524 4238 20580
rect 4498 20524 4508 20580
rect 4564 20524 6300 20580
rect 6356 20524 6366 20580
rect 8530 20524 8540 20580
rect 8596 20524 9436 20580
rect 9492 20524 9502 20580
rect 18610 20524 18620 20580
rect 18676 20524 20636 20580
rect 20692 20524 21196 20580
rect 21252 20524 21262 20580
rect 31826 20524 31836 20580
rect 31892 20524 33292 20580
rect 33348 20524 33358 20580
rect 34486 20524 34524 20580
rect 34580 20524 34590 20580
rect 5842 20412 5852 20468
rect 5908 20412 11340 20468
rect 11396 20412 12236 20468
rect 12292 20412 13468 20468
rect 13524 20412 13534 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 2940 20300 4844 20356
rect 4900 20300 5348 20356
rect 9538 20300 9548 20356
rect 9604 20300 10556 20356
rect 10612 20300 10622 20356
rect 33842 20300 33852 20356
rect 33908 20300 34188 20356
rect 34244 20300 34254 20356
rect 0 20244 800 20272
rect 0 20188 1708 20244
rect 1764 20188 2492 20244
rect 2548 20188 2558 20244
rect 0 20160 800 20188
rect 2940 20132 2996 20300
rect 3154 20188 3164 20244
rect 3220 20188 3836 20244
rect 3892 20188 3902 20244
rect 5292 20132 5348 20300
rect 41101 20244 41901 20272
rect 13794 20188 13804 20244
rect 13860 20188 13870 20244
rect 18162 20188 18172 20244
rect 18228 20188 18238 20244
rect 20738 20188 20748 20244
rect 20804 20188 21644 20244
rect 21700 20188 21710 20244
rect 31836 20188 36428 20244
rect 36484 20188 37212 20244
rect 37268 20188 37278 20244
rect 39676 20188 41901 20244
rect 13804 20132 13860 20188
rect 18172 20132 18228 20188
rect 31836 20132 31892 20188
rect 39676 20132 39732 20188
rect 41101 20160 41901 20188
rect 2940 20076 3276 20132
rect 3332 20076 3342 20132
rect 3714 20076 3724 20132
rect 3780 20076 3790 20132
rect 5282 20076 5292 20132
rect 5348 20076 5358 20132
rect 10882 20076 10892 20132
rect 10948 20076 10958 20132
rect 13122 20076 13132 20132
rect 13188 20076 14588 20132
rect 14644 20076 14654 20132
rect 18060 20076 18228 20132
rect 18946 20076 18956 20132
rect 19012 20076 19292 20132
rect 19348 20076 19740 20132
rect 19796 20076 20412 20132
rect 20468 20076 20478 20132
rect 20962 20076 20972 20132
rect 21028 20076 21756 20132
rect 21812 20076 21822 20132
rect 29362 20076 29372 20132
rect 29428 20076 31892 20132
rect 33394 20076 33404 20132
rect 33460 20076 38892 20132
rect 38948 20076 38958 20132
rect 39666 20076 39676 20132
rect 39732 20076 39742 20132
rect 3724 20020 3780 20076
rect 10892 20020 10948 20076
rect 2706 19964 2716 20020
rect 2772 19964 3780 20020
rect 4050 19964 4060 20020
rect 4116 19964 4956 20020
rect 5012 19964 6188 20020
rect 6244 19964 6254 20020
rect 8194 19964 8204 20020
rect 8260 19964 8652 20020
rect 8708 19964 9324 20020
rect 9380 19964 10948 20020
rect 11106 19964 11116 20020
rect 11172 19964 12236 20020
rect 12292 19964 12302 20020
rect 12562 19964 12572 20020
rect 12628 19964 14252 20020
rect 14308 19964 14318 20020
rect 3042 19852 3052 19908
rect 3108 19852 3388 19908
rect 4722 19852 4732 19908
rect 4788 19852 5292 19908
rect 5348 19852 5358 19908
rect 8390 19852 8428 19908
rect 8484 19852 8494 19908
rect 8978 19852 8988 19908
rect 9044 19852 9436 19908
rect 9492 19852 9660 19908
rect 9716 19852 9726 19908
rect 12114 19852 12124 19908
rect 12180 19852 13356 19908
rect 13412 19852 14476 19908
rect 14532 19852 14542 19908
rect 0 19572 800 19600
rect 0 19516 1708 19572
rect 1764 19516 2492 19572
rect 2548 19516 2558 19572
rect 0 19488 800 19516
rect 3332 19460 3388 19852
rect 18060 19796 18116 20076
rect 18274 19964 18284 20020
rect 18340 19964 20860 20020
rect 20916 19964 20926 20020
rect 26674 19964 26684 20020
rect 26740 19964 27020 20020
rect 27076 19964 27086 20020
rect 27234 19964 27244 20020
rect 27300 19964 27310 20020
rect 28354 19964 28364 20020
rect 28420 19964 29932 20020
rect 29988 19964 30380 20020
rect 30436 19964 30446 20020
rect 31378 19964 31388 20020
rect 31444 19964 32508 20020
rect 32564 19964 32956 20020
rect 33012 19964 33516 20020
rect 33572 19964 33582 20020
rect 33730 19964 33740 20020
rect 33796 19964 34860 20020
rect 34916 19964 34926 20020
rect 35410 19964 35420 20020
rect 35476 19964 36876 20020
rect 36932 19964 36942 20020
rect 27244 19908 27300 19964
rect 19058 19852 19068 19908
rect 19124 19852 19628 19908
rect 19684 19852 19694 19908
rect 25218 19852 25228 19908
rect 25284 19852 25900 19908
rect 25956 19852 25966 19908
rect 26450 19852 26460 19908
rect 26516 19852 27300 19908
rect 27458 19852 27468 19908
rect 27524 19852 38668 19908
rect 38612 19796 38668 19852
rect 18022 19740 18060 19796
rect 18116 19740 26348 19796
rect 26404 19740 26414 19796
rect 26852 19740 28140 19796
rect 28196 19740 31724 19796
rect 31780 19740 31790 19796
rect 33814 19740 33852 19796
rect 33908 19740 33918 19796
rect 34514 19740 34524 19796
rect 34580 19740 34590 19796
rect 38612 19740 39116 19796
rect 39172 19740 39182 19796
rect 9314 19628 9324 19684
rect 9380 19628 13580 19684
rect 13636 19628 13646 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 26852 19572 26908 19740
rect 34524 19684 34580 19740
rect 27010 19628 27020 19684
rect 27076 19628 34580 19684
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41101 19572 41901 19600
rect 24658 19516 24668 19572
rect 24724 19516 26908 19572
rect 28690 19516 28700 19572
rect 28756 19516 29484 19572
rect 29540 19516 31276 19572
rect 31332 19516 31342 19572
rect 40002 19516 40012 19572
rect 40068 19516 41901 19572
rect 41101 19488 41901 19516
rect 3332 19404 4620 19460
rect 4676 19404 6524 19460
rect 6580 19404 6590 19460
rect 12786 19404 12796 19460
rect 12852 19404 13468 19460
rect 13524 19404 13534 19460
rect 21634 19404 21644 19460
rect 21700 19404 23772 19460
rect 23828 19404 26236 19460
rect 26292 19404 26302 19460
rect 26562 19404 26572 19460
rect 26628 19404 29260 19460
rect 29316 19404 29326 19460
rect 2818 19292 2828 19348
rect 2884 19292 3388 19348
rect 4722 19292 4732 19348
rect 4788 19292 4844 19348
rect 4900 19292 4910 19348
rect 14028 19292 17388 19348
rect 17444 19292 17454 19348
rect 3332 18676 3388 19292
rect 14028 19236 14084 19292
rect 8306 19180 8316 19236
rect 8372 19180 8988 19236
rect 9044 19180 9054 19236
rect 9426 19180 9436 19236
rect 9492 19180 9884 19236
rect 9940 19180 12572 19236
rect 12628 19180 12638 19236
rect 14018 19180 14028 19236
rect 14084 19180 14094 19236
rect 15362 19180 15372 19236
rect 15428 19180 23660 19236
rect 23716 19180 24332 19236
rect 24388 19180 24398 19236
rect 25218 19180 25228 19236
rect 25284 19180 28588 19236
rect 28644 19180 29260 19236
rect 29316 19180 29326 19236
rect 36530 19180 36540 19236
rect 36596 19180 37436 19236
rect 37492 19180 37502 19236
rect 6402 19068 6412 19124
rect 6468 19068 7532 19124
rect 7588 19068 7598 19124
rect 8418 19068 8428 19124
rect 8484 19068 9660 19124
rect 9716 19068 9726 19124
rect 19590 19068 19628 19124
rect 19684 19068 19964 19124
rect 20020 19068 20030 19124
rect 30594 19068 30604 19124
rect 30660 19068 31276 19124
rect 31332 19068 31342 19124
rect 32946 19068 32956 19124
rect 33012 19068 34412 19124
rect 34468 19068 34478 19124
rect 3602 18956 3612 19012
rect 3668 18956 6300 19012
rect 6356 18956 6366 19012
rect 6626 18956 6636 19012
rect 6692 18956 7420 19012
rect 7476 18956 7486 19012
rect 7746 18956 7756 19012
rect 7812 18956 8428 19012
rect 8484 18956 8494 19012
rect 17378 18956 17388 19012
rect 17444 18956 17836 19012
rect 17892 18956 17902 19012
rect 18946 18956 18956 19012
rect 19012 18956 19180 19012
rect 19236 18956 19246 19012
rect 19394 18956 19404 19012
rect 19460 18956 20300 19012
rect 20356 18956 20366 19012
rect 6076 18900 6132 18956
rect 41101 18900 41901 18928
rect 6066 18844 6076 18900
rect 6132 18844 6142 18900
rect 8642 18844 8652 18900
rect 8708 18844 8988 18900
rect 9044 18844 18956 18900
rect 19012 18844 19022 18900
rect 20178 18844 20188 18900
rect 20244 18844 21028 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 5394 18732 5404 18788
rect 5460 18732 6412 18788
rect 6468 18732 6478 18788
rect 20188 18676 20244 18844
rect 20972 18676 21028 18844
rect 26852 18844 33628 18900
rect 33684 18844 33694 18900
rect 39666 18844 39676 18900
rect 39732 18844 41901 18900
rect 26852 18676 26908 18844
rect 41101 18816 41901 18844
rect 3332 18620 10108 18676
rect 10164 18620 10174 18676
rect 18834 18620 18844 18676
rect 18900 18620 20244 18676
rect 20962 18620 20972 18676
rect 21028 18620 26908 18676
rect 29810 18620 29820 18676
rect 29876 18620 37324 18676
rect 37380 18620 37390 18676
rect 4172 18452 4228 18620
rect 6262 18508 6300 18564
rect 6356 18508 6366 18564
rect 7634 18508 7644 18564
rect 7700 18508 8428 18564
rect 8484 18508 9436 18564
rect 9492 18508 9502 18564
rect 18498 18508 18508 18564
rect 18564 18508 19740 18564
rect 19796 18508 20412 18564
rect 20468 18508 20478 18564
rect 33730 18508 33740 18564
rect 33796 18508 34636 18564
rect 34692 18508 34702 18564
rect 36642 18508 36652 18564
rect 36708 18508 37772 18564
rect 37828 18508 37838 18564
rect 1922 18396 1932 18452
rect 1988 18396 3724 18452
rect 3780 18396 3790 18452
rect 4162 18396 4172 18452
rect 4228 18396 4238 18452
rect 7186 18396 7196 18452
rect 7252 18396 8204 18452
rect 8260 18396 8270 18452
rect 10322 18396 10332 18452
rect 10388 18396 12796 18452
rect 12852 18396 12862 18452
rect 13010 18396 13020 18452
rect 13076 18396 13692 18452
rect 13748 18396 13758 18452
rect 17042 18396 17052 18452
rect 17108 18396 17836 18452
rect 17892 18396 20524 18452
rect 20580 18396 20590 18452
rect 24770 18396 24780 18452
rect 24836 18396 25340 18452
rect 25396 18396 25406 18452
rect 26674 18396 26684 18452
rect 26740 18396 27244 18452
rect 27300 18396 27310 18452
rect 32498 18396 32508 18452
rect 32564 18396 34300 18452
rect 34356 18396 34366 18452
rect 36978 18396 36988 18452
rect 37044 18396 37996 18452
rect 38052 18396 38062 18452
rect 38612 18396 38892 18452
rect 38948 18396 38958 18452
rect 38612 18340 38668 18396
rect 12226 18284 12236 18340
rect 12292 18284 13244 18340
rect 13300 18284 17388 18340
rect 17444 18284 17612 18340
rect 17668 18284 17678 18340
rect 25106 18284 25116 18340
rect 25172 18284 25564 18340
rect 25620 18284 25630 18340
rect 34850 18284 34860 18340
rect 34916 18284 36316 18340
rect 36372 18284 36382 18340
rect 37426 18284 37436 18340
rect 37492 18284 38668 18340
rect 41101 18228 41901 18256
rect 4498 18172 4508 18228
rect 4564 18172 5404 18228
rect 5460 18172 5470 18228
rect 6860 18172 7532 18228
rect 7588 18172 8204 18228
rect 8260 18172 8270 18228
rect 14242 18172 14252 18228
rect 14308 18172 24892 18228
rect 24948 18172 24958 18228
rect 34066 18172 34076 18228
rect 34132 18172 34636 18228
rect 34692 18172 35308 18228
rect 35364 18172 35374 18228
rect 38098 18172 38108 18228
rect 38164 18172 41901 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 6860 18004 6916 18172
rect 41101 18144 41901 18172
rect 12898 18060 12908 18116
rect 12964 18060 19404 18116
rect 19460 18060 23884 18116
rect 23940 18060 24332 18116
rect 24388 18060 24398 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 6178 17948 6188 18004
rect 6244 17948 6860 18004
rect 6916 17948 6926 18004
rect 16818 17948 16828 18004
rect 16884 17948 18620 18004
rect 18676 17948 19292 18004
rect 19348 17948 19358 18004
rect 17798 17836 17836 17892
rect 17892 17836 17902 17892
rect 19058 17836 19068 17892
rect 19124 17836 19628 17892
rect 19684 17836 19694 17892
rect 34514 17836 34524 17892
rect 34580 17836 36092 17892
rect 36148 17836 36158 17892
rect 21522 17724 21532 17780
rect 21588 17724 24556 17780
rect 24612 17724 25228 17780
rect 25284 17724 25564 17780
rect 25620 17724 25630 17780
rect 28924 17724 38556 17780
rect 38612 17724 38622 17780
rect 14466 17612 14476 17668
rect 14532 17612 16044 17668
rect 16100 17612 16110 17668
rect 28924 17556 28980 17724
rect 29138 17612 29148 17668
rect 29204 17612 29484 17668
rect 29540 17612 31500 17668
rect 31556 17612 31566 17668
rect 41101 17556 41901 17584
rect 27122 17500 27132 17556
rect 27188 17500 28980 17556
rect 30482 17500 30492 17556
rect 30548 17500 31164 17556
rect 31220 17500 31230 17556
rect 33058 17500 33068 17556
rect 33124 17500 33852 17556
rect 33908 17500 33918 17556
rect 39666 17500 39676 17556
rect 39732 17500 41901 17556
rect 41101 17472 41901 17500
rect 15474 17388 15484 17444
rect 15540 17388 16716 17444
rect 16772 17388 16782 17444
rect 23202 17388 23212 17444
rect 23268 17388 26684 17444
rect 26740 17388 30716 17444
rect 30772 17388 30782 17444
rect 32162 17388 32172 17444
rect 32228 17388 35084 17444
rect 35140 17388 35150 17444
rect 34290 17276 34300 17332
rect 34356 17276 40012 17332
rect 40068 17276 40078 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 5618 17164 5628 17220
rect 5684 17164 5964 17220
rect 6020 17164 6030 17220
rect 33394 17052 33404 17108
rect 33460 17052 33852 17108
rect 33908 17052 34972 17108
rect 35028 17052 35038 17108
rect 35970 17052 35980 17108
rect 36036 17052 36764 17108
rect 36820 17052 36830 17108
rect 28466 16940 28476 16996
rect 28532 16940 29148 16996
rect 29204 16940 29214 16996
rect 29922 16940 29932 16996
rect 29988 16940 30492 16996
rect 30548 16940 30558 16996
rect 31938 16940 31948 16996
rect 32004 16940 32014 16996
rect 34626 16940 34636 16996
rect 34692 16940 35812 16996
rect 36642 16940 36652 16996
rect 36708 16940 37996 16996
rect 38052 16940 38062 16996
rect 7494 16828 7532 16884
rect 7588 16828 7598 16884
rect 7746 16828 7756 16884
rect 7812 16828 8764 16884
rect 8820 16828 8830 16884
rect 31948 16772 32004 16940
rect 34738 16828 34748 16884
rect 34804 16828 35532 16884
rect 35588 16828 35598 16884
rect 35756 16772 35812 16940
rect 41101 16884 41901 16912
rect 36194 16828 36204 16884
rect 36260 16828 37212 16884
rect 37268 16828 37278 16884
rect 39778 16828 39788 16884
rect 39844 16828 41901 16884
rect 41101 16800 41901 16828
rect 16706 16716 16716 16772
rect 16772 16716 17052 16772
rect 17108 16716 19068 16772
rect 19124 16716 19134 16772
rect 31948 16716 32844 16772
rect 32900 16716 32910 16772
rect 33506 16716 33516 16772
rect 33572 16716 34188 16772
rect 34244 16716 35196 16772
rect 35252 16716 35262 16772
rect 35756 16716 38668 16772
rect 3602 16604 3612 16660
rect 3668 16604 7532 16660
rect 7588 16604 7598 16660
rect 38612 16548 38668 16716
rect 4946 16492 4956 16548
rect 5012 16492 5628 16548
rect 5684 16492 5852 16548
rect 5908 16492 6748 16548
rect 6804 16492 6814 16548
rect 18498 16492 18508 16548
rect 18564 16492 18788 16548
rect 38612 16492 40124 16548
rect 40180 16492 40190 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 4834 16380 4844 16436
rect 4900 16380 5740 16436
rect 5796 16380 11564 16436
rect 11620 16380 11630 16436
rect 4610 16268 4620 16324
rect 4676 16268 6188 16324
rect 6244 16268 6254 16324
rect 16818 16268 16828 16324
rect 16884 16268 17948 16324
rect 18004 16268 18508 16324
rect 18564 16268 18574 16324
rect 18732 16212 18788 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 27906 16268 27916 16324
rect 27972 16268 28588 16324
rect 28644 16268 28654 16324
rect 35074 16268 35084 16324
rect 35140 16268 38892 16324
rect 38948 16268 38958 16324
rect 41101 16212 41901 16240
rect 6290 16156 6300 16212
rect 6356 16156 7308 16212
rect 7364 16156 7374 16212
rect 8082 16156 8092 16212
rect 8148 16156 8540 16212
rect 8596 16156 8606 16212
rect 18722 16156 18732 16212
rect 18788 16156 18798 16212
rect 22306 16156 22316 16212
rect 22372 16156 22876 16212
rect 22932 16156 25004 16212
rect 25060 16156 25070 16212
rect 30146 16156 30156 16212
rect 30212 16156 37436 16212
rect 37492 16156 37502 16212
rect 38322 16156 38332 16212
rect 38388 16156 41901 16212
rect 41101 16128 41901 16156
rect 6402 16044 6412 16100
rect 6468 16044 7084 16100
rect 7140 16044 7150 16100
rect 19506 16044 19516 16100
rect 19572 16044 25116 16100
rect 25172 16044 25676 16100
rect 25732 16044 25742 16100
rect 30818 16044 30828 16100
rect 30884 16044 37324 16100
rect 37380 16044 37390 16100
rect 6962 15932 6972 15988
rect 7028 15932 7644 15988
rect 7700 15932 7710 15988
rect 20066 15932 20076 15988
rect 20132 15932 23436 15988
rect 23492 15932 24332 15988
rect 24388 15932 24780 15988
rect 24836 15932 24846 15988
rect 31938 15932 31948 15988
rect 32004 15932 33068 15988
rect 33124 15932 33134 15988
rect 17602 15820 17612 15876
rect 17668 15820 18060 15876
rect 18116 15820 18126 15876
rect 19254 15820 19292 15876
rect 19348 15820 19358 15876
rect 29474 15820 29484 15876
rect 29540 15820 37324 15876
rect 37380 15820 37390 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 23090 15596 23100 15652
rect 23156 15596 33292 15652
rect 33348 15596 34300 15652
rect 34356 15596 34366 15652
rect 41101 15540 41901 15568
rect 5954 15484 5964 15540
rect 6020 15484 6030 15540
rect 7746 15484 7756 15540
rect 7812 15484 8316 15540
rect 8372 15484 8382 15540
rect 9090 15484 9100 15540
rect 9156 15484 9772 15540
rect 9828 15484 9838 15540
rect 12450 15484 12460 15540
rect 12516 15484 13916 15540
rect 13972 15484 16044 15540
rect 16100 15484 16110 15540
rect 16370 15484 16380 15540
rect 16436 15484 16604 15540
rect 16660 15484 16670 15540
rect 19730 15484 19740 15540
rect 19796 15484 22092 15540
rect 22148 15484 22158 15540
rect 32834 15484 32844 15540
rect 32900 15484 38892 15540
rect 38948 15484 38958 15540
rect 39554 15484 39564 15540
rect 39620 15484 41901 15540
rect 5964 15316 6020 15484
rect 41101 15456 41901 15484
rect 7074 15372 7084 15428
rect 7140 15372 7644 15428
rect 7700 15372 8204 15428
rect 8260 15372 8270 15428
rect 8418 15372 8428 15428
rect 8484 15372 8522 15428
rect 16706 15372 16716 15428
rect 16772 15372 18172 15428
rect 18228 15372 18396 15428
rect 18452 15372 18462 15428
rect 5506 15260 5516 15316
rect 5572 15260 7868 15316
rect 7924 15260 7934 15316
rect 8754 15260 8764 15316
rect 8820 15260 9772 15316
rect 9828 15260 9838 15316
rect 19058 15260 19068 15316
rect 19124 15260 19628 15316
rect 19684 15260 19694 15316
rect 31042 15260 31052 15316
rect 31108 15260 31388 15316
rect 31444 15260 32172 15316
rect 32228 15260 32238 15316
rect 6962 15148 6972 15204
rect 7028 15148 7196 15204
rect 7252 15148 11900 15204
rect 11956 15148 11966 15204
rect 23874 15148 23884 15204
rect 23940 15148 25340 15204
rect 25396 15148 25406 15204
rect 30034 15148 30044 15204
rect 30100 15148 31332 15204
rect 31276 15092 31332 15148
rect 12450 15036 12460 15092
rect 12516 15036 14364 15092
rect 14420 15036 14430 15092
rect 18050 15036 18060 15092
rect 18116 15036 29932 15092
rect 29988 15036 29998 15092
rect 30146 15036 30156 15092
rect 30212 15036 31052 15092
rect 31108 15036 31118 15092
rect 31276 15036 38892 15092
rect 38948 15036 38958 15092
rect 17378 14924 17388 14980
rect 17444 14924 18508 14980
rect 18564 14924 18574 14980
rect 18946 14924 18956 14980
rect 19012 14924 19964 14980
rect 20020 14924 20030 14980
rect 31154 14924 31164 14980
rect 31220 14924 31612 14980
rect 31668 14924 31678 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 41101 14868 41901 14896
rect 15026 14812 15036 14868
rect 15092 14812 15372 14868
rect 15428 14812 18396 14868
rect 18452 14812 18462 14868
rect 20738 14812 20748 14868
rect 20804 14812 21420 14868
rect 21476 14812 28700 14868
rect 28756 14812 28766 14868
rect 30482 14812 30492 14868
rect 30548 14812 30940 14868
rect 30996 14812 31006 14868
rect 38098 14812 38108 14868
rect 38164 14812 41901 14868
rect 41101 14784 41901 14812
rect 9398 14700 9436 14756
rect 9492 14700 9502 14756
rect 17938 14700 17948 14756
rect 18004 14700 18956 14756
rect 19012 14700 19022 14756
rect 29810 14700 29820 14756
rect 29876 14700 32060 14756
rect 32116 14700 33404 14756
rect 33460 14700 33470 14756
rect 5058 14588 5068 14644
rect 5124 14588 5516 14644
rect 5572 14588 5852 14644
rect 5908 14588 5918 14644
rect 27234 14588 27244 14644
rect 27300 14588 29148 14644
rect 29204 14588 29214 14644
rect 4834 14476 4844 14532
rect 4900 14476 5964 14532
rect 6020 14476 6972 14532
rect 7028 14476 7038 14532
rect 12338 14476 12348 14532
rect 12404 14476 14028 14532
rect 14084 14476 14094 14532
rect 22754 14476 22764 14532
rect 22820 14476 23324 14532
rect 23380 14476 23772 14532
rect 23828 14476 23838 14532
rect 23986 14476 23996 14532
rect 24052 14476 25116 14532
rect 25172 14476 27132 14532
rect 27188 14476 27198 14532
rect 6626 14364 6636 14420
rect 6692 14364 8428 14420
rect 8484 14364 8494 14420
rect 13458 14364 13468 14420
rect 13524 14364 15372 14420
rect 15428 14364 15438 14420
rect 16146 14364 16156 14420
rect 16212 14364 17948 14420
rect 18004 14364 18014 14420
rect 19282 14364 19292 14420
rect 19348 14364 19740 14420
rect 19796 14364 19806 14420
rect 12898 14252 12908 14308
rect 12964 14252 13692 14308
rect 13748 14252 16716 14308
rect 16772 14252 17500 14308
rect 17556 14252 17566 14308
rect 18386 14252 18396 14308
rect 18452 14252 20356 14308
rect 25890 14252 25900 14308
rect 25956 14252 26796 14308
rect 26852 14252 26862 14308
rect 20300 14196 20356 14252
rect 20300 14140 20748 14196
rect 20804 14140 20814 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 20300 14084 20356 14140
rect 3332 14028 8540 14084
rect 8596 14028 8606 14084
rect 20290 14028 20300 14084
rect 20356 14028 20366 14084
rect 23426 14028 23436 14084
rect 23492 14028 25340 14084
rect 25396 14028 25406 14084
rect 32162 14028 32172 14084
rect 32228 14028 33516 14084
rect 33572 14028 33582 14084
rect 3332 13860 3388 14028
rect 8642 13916 8652 13972
rect 8708 13916 9212 13972
rect 9268 13916 9660 13972
rect 9716 13916 9726 13972
rect 13458 13916 13468 13972
rect 13524 13916 15596 13972
rect 15652 13916 15662 13972
rect 18274 13916 18284 13972
rect 18340 13916 19068 13972
rect 19124 13916 19134 13972
rect 20738 13916 20748 13972
rect 20804 13916 22204 13972
rect 22260 13916 22270 13972
rect 24658 13916 24668 13972
rect 24724 13916 25452 13972
rect 25508 13916 25518 13972
rect 28802 13916 28812 13972
rect 28868 13916 29820 13972
rect 29876 13916 30156 13972
rect 30212 13916 30222 13972
rect 20748 13860 20804 13916
rect 2482 13804 2492 13860
rect 2548 13804 3388 13860
rect 8194 13804 8204 13860
rect 8260 13804 9996 13860
rect 10052 13804 10062 13860
rect 14028 13804 17388 13860
rect 17444 13804 17454 13860
rect 17826 13804 17836 13860
rect 17892 13804 19180 13860
rect 19236 13804 20804 13860
rect 30370 13804 30380 13860
rect 30436 13804 30446 13860
rect 33058 13804 33068 13860
rect 33124 13804 33134 13860
rect 34626 13804 34636 13860
rect 34692 13804 35644 13860
rect 35700 13804 35710 13860
rect 14028 13748 14084 13804
rect 9286 13692 9324 13748
rect 9380 13692 9390 13748
rect 11442 13692 11452 13748
rect 11508 13692 12460 13748
rect 12516 13692 12526 13748
rect 13346 13692 13356 13748
rect 13412 13692 14028 13748
rect 14084 13692 14094 13748
rect 14914 13692 14924 13748
rect 14980 13692 15932 13748
rect 15988 13692 16828 13748
rect 16884 13692 17612 13748
rect 17668 13692 17678 13748
rect 10322 13580 10332 13636
rect 10388 13580 11004 13636
rect 11060 13580 13804 13636
rect 13860 13580 13870 13636
rect 14690 13580 14700 13636
rect 14756 13580 15484 13636
rect 15540 13580 15550 13636
rect 17948 13580 18956 13636
rect 19012 13580 19022 13636
rect 26674 13580 26684 13636
rect 26740 13580 28252 13636
rect 28308 13580 28318 13636
rect 17948 13524 18004 13580
rect 11330 13468 11340 13524
rect 11396 13468 12012 13524
rect 12068 13468 12078 13524
rect 14242 13468 14252 13524
rect 14308 13468 15036 13524
rect 15092 13468 18004 13524
rect 18162 13468 18172 13524
rect 18228 13468 19516 13524
rect 19572 13468 19582 13524
rect 26002 13468 26012 13524
rect 26068 13468 27468 13524
rect 27524 13468 27534 13524
rect 30380 13412 30436 13804
rect 33068 13636 33124 13804
rect 32050 13580 32060 13636
rect 32116 13580 33124 13636
rect 30706 13468 30716 13524
rect 30772 13468 31612 13524
rect 31668 13468 31678 13524
rect 8082 13356 8092 13412
rect 8148 13356 8540 13412
rect 8596 13356 8606 13412
rect 17154 13356 17164 13412
rect 17220 13356 18060 13412
rect 18116 13356 18126 13412
rect 21298 13356 21308 13412
rect 21364 13356 21374 13412
rect 21858 13356 21868 13412
rect 21924 13356 30436 13412
rect 30594 13356 30604 13412
rect 30660 13356 31388 13412
rect 31444 13356 31454 13412
rect 31892 13356 32508 13412
rect 32564 13356 32574 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 21308 13300 21364 13356
rect 31892 13300 31948 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 17938 13244 17948 13300
rect 18004 13244 21364 13300
rect 28914 13244 28924 13300
rect 28980 13244 31948 13300
rect 7410 13132 7420 13188
rect 7476 13132 9660 13188
rect 9716 13132 9726 13188
rect 25218 13132 25228 13188
rect 25284 13132 27244 13188
rect 27300 13132 27916 13188
rect 27972 13132 27982 13188
rect 5842 13020 5852 13076
rect 5908 13020 6188 13076
rect 6244 13020 7644 13076
rect 7700 13020 7710 13076
rect 4834 12908 4844 12964
rect 4900 12908 5516 12964
rect 5572 12908 5582 12964
rect 16706 12908 16716 12964
rect 16772 12908 21196 12964
rect 21252 12908 21262 12964
rect 30828 12852 30884 13244
rect 32162 13132 32172 13188
rect 32228 13132 33068 13188
rect 33124 13132 33292 13188
rect 33348 13132 33964 13188
rect 34020 13132 34030 13188
rect 31266 13020 31276 13076
rect 31332 13020 38948 13076
rect 38892 12964 38948 13020
rect 31042 12908 31052 12964
rect 31108 12908 32620 12964
rect 32676 12908 32686 12964
rect 38882 12908 38892 12964
rect 38948 12908 38958 12964
rect 41101 12852 41901 12880
rect 9538 12796 9548 12852
rect 9604 12796 10444 12852
rect 10500 12796 10510 12852
rect 30828 12796 31164 12852
rect 31220 12796 31230 12852
rect 34066 12796 34076 12852
rect 34132 12796 35644 12852
rect 35700 12796 35710 12852
rect 40002 12796 40012 12852
rect 40068 12796 41901 12852
rect 41101 12768 41901 12796
rect 7970 12684 7980 12740
rect 8036 12684 8988 12740
rect 9044 12684 9054 12740
rect 11890 12684 11900 12740
rect 11956 12684 13580 12740
rect 13636 12684 13646 12740
rect 36418 12684 36428 12740
rect 36484 12684 37100 12740
rect 37156 12684 37166 12740
rect 9874 12572 9884 12628
rect 9940 12572 11564 12628
rect 11620 12572 12572 12628
rect 12628 12572 12638 12628
rect 19170 12572 19180 12628
rect 19236 12572 19516 12628
rect 19572 12572 19582 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 12226 12460 12236 12516
rect 12292 12460 13468 12516
rect 13524 12460 13534 12516
rect 15586 12460 15596 12516
rect 15652 12460 15662 12516
rect 6626 12348 6636 12404
rect 6692 12348 8764 12404
rect 8820 12348 9996 12404
rect 10052 12348 11788 12404
rect 11844 12348 11854 12404
rect 13570 12348 13580 12404
rect 13636 12348 15260 12404
rect 15316 12348 15326 12404
rect 15596 12292 15652 12460
rect 18946 12348 18956 12404
rect 19012 12348 23212 12404
rect 23268 12348 23278 12404
rect 4834 12236 4844 12292
rect 4900 12236 6076 12292
rect 6132 12236 6142 12292
rect 14018 12236 14028 12292
rect 14084 12236 15652 12292
rect 19730 12236 19740 12292
rect 19796 12236 20300 12292
rect 20356 12236 20636 12292
rect 20692 12236 20702 12292
rect 41101 12180 41901 12208
rect 5730 12124 5740 12180
rect 5796 12124 7756 12180
rect 7812 12124 7822 12180
rect 14130 12124 14140 12180
rect 14196 12124 15708 12180
rect 15764 12124 15774 12180
rect 17826 12124 17836 12180
rect 17892 12124 19404 12180
rect 19460 12124 19470 12180
rect 28018 12124 28028 12180
rect 28084 12124 28588 12180
rect 28644 12124 29820 12180
rect 29876 12124 31612 12180
rect 31668 12124 33516 12180
rect 33572 12124 33582 12180
rect 40114 12124 40124 12180
rect 40180 12124 41901 12180
rect 41101 12096 41901 12124
rect 4498 12012 4508 12068
rect 4564 12012 4956 12068
rect 5012 12012 5022 12068
rect 8082 12012 8092 12068
rect 8148 12012 9660 12068
rect 9716 12012 9726 12068
rect 13122 12012 13132 12068
rect 13188 12012 14588 12068
rect 14644 12012 15148 12068
rect 15204 12012 15214 12068
rect 16594 12012 16604 12068
rect 16660 12012 18508 12068
rect 18564 12012 19292 12068
rect 19348 12012 19358 12068
rect 6738 11900 6748 11956
rect 6804 11900 10668 11956
rect 10724 11900 14028 11956
rect 14084 11900 14094 11956
rect 24322 11900 24332 11956
rect 24388 11900 25228 11956
rect 25284 11900 25294 11956
rect 25554 11900 25564 11956
rect 25620 11900 26348 11956
rect 26404 11900 26414 11956
rect 15698 11788 15708 11844
rect 15764 11788 17836 11844
rect 17892 11788 18732 11844
rect 18788 11788 24444 11844
rect 24500 11788 24510 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 5842 11676 5852 11732
rect 5908 11676 7196 11732
rect 7252 11676 11228 11732
rect 11284 11676 11294 11732
rect 14018 11676 14028 11732
rect 14084 11676 16156 11732
rect 16212 11676 16222 11732
rect 16930 11676 16940 11732
rect 16996 11676 18172 11732
rect 18228 11676 18238 11732
rect 16482 11564 16492 11620
rect 16548 11564 17612 11620
rect 17668 11564 17678 11620
rect 9426 11452 9436 11508
rect 9492 11452 10556 11508
rect 10612 11452 11900 11508
rect 11956 11452 11966 11508
rect 15138 11452 15148 11508
rect 15204 11452 20188 11508
rect 20244 11452 20524 11508
rect 20580 11452 21084 11508
rect 21140 11452 21150 11508
rect 7522 11340 7532 11396
rect 7588 11340 8428 11396
rect 8484 11340 8494 11396
rect 8754 11340 8764 11396
rect 8820 11340 9212 11396
rect 9268 11340 11172 11396
rect 12898 11340 12908 11396
rect 12964 11340 13580 11396
rect 13636 11340 13646 11396
rect 16818 11340 16828 11396
rect 16884 11340 17836 11396
rect 17892 11340 17902 11396
rect 24994 11340 25004 11396
rect 25060 11340 30940 11396
rect 30996 11340 32956 11396
rect 33012 11340 33516 11396
rect 33572 11340 33582 11396
rect 11116 11284 11172 11340
rect 5954 11228 5964 11284
rect 6020 11228 6748 11284
rect 6804 11228 6814 11284
rect 9090 11228 9100 11284
rect 9156 11228 10108 11284
rect 10164 11228 10174 11284
rect 11116 11228 14588 11284
rect 14644 11228 14654 11284
rect 16930 11228 16940 11284
rect 16996 11228 17948 11284
rect 18004 11228 20076 11284
rect 20132 11228 21308 11284
rect 21364 11228 21374 11284
rect 28242 11228 28252 11284
rect 28308 11228 29484 11284
rect 29540 11228 30044 11284
rect 30100 11228 30110 11284
rect 31714 11228 31724 11284
rect 31780 11228 32844 11284
rect 32900 11228 33292 11284
rect 33348 11228 33358 11284
rect 8754 11116 8764 11172
rect 8820 11116 9772 11172
rect 9828 11116 9838 11172
rect 16034 11116 16044 11172
rect 16100 11116 17388 11172
rect 17444 11116 17454 11172
rect 27906 11116 27916 11172
rect 27972 11116 28588 11172
rect 28644 11116 28654 11172
rect 30818 11116 30828 11172
rect 30884 11116 31388 11172
rect 31444 11116 31836 11172
rect 31892 11116 31902 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 3332 10892 8372 10948
rect 3332 10836 3388 10892
rect 8316 10836 8372 10892
rect 2706 10780 2716 10836
rect 2772 10780 3388 10836
rect 4946 10780 4956 10836
rect 5012 10780 6300 10836
rect 6356 10780 6366 10836
rect 8306 10780 8316 10836
rect 8372 10780 8382 10836
rect 9986 10668 9996 10724
rect 10052 10668 10556 10724
rect 10612 10668 17052 10724
rect 17108 10668 19964 10724
rect 20020 10668 20030 10724
rect 28242 10668 28252 10724
rect 28308 10668 28924 10724
rect 28980 10668 29708 10724
rect 29764 10668 29774 10724
rect 3042 10556 3052 10612
rect 3108 10556 10108 10612
rect 10164 10556 10174 10612
rect 10322 10556 10332 10612
rect 10388 10556 12124 10612
rect 12180 10556 12190 10612
rect 24546 10556 24556 10612
rect 24612 10556 25340 10612
rect 25396 10556 25406 10612
rect 29474 10556 29484 10612
rect 29540 10556 30268 10612
rect 30324 10556 30334 10612
rect 2370 10444 2380 10500
rect 2436 10444 4956 10500
rect 5012 10444 5022 10500
rect 8194 10444 8204 10500
rect 8260 10444 8876 10500
rect 8932 10444 8942 10500
rect 34066 10444 34076 10500
rect 34132 10444 35644 10500
rect 35700 10444 35710 10500
rect 31714 10332 31724 10388
rect 31780 10332 32732 10388
rect 32788 10332 32798 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 20402 10108 20412 10164
rect 20468 10108 21420 10164
rect 21476 10108 21868 10164
rect 21924 10108 23660 10164
rect 23716 10108 23726 10164
rect 19282 9996 19292 10052
rect 19348 9996 19740 10052
rect 19796 9996 26236 10052
rect 26292 9996 26302 10052
rect 20738 9884 20748 9940
rect 20804 9884 21532 9940
rect 21588 9884 23436 9940
rect 23492 9884 23502 9940
rect 23650 9884 23660 9940
rect 23716 9884 25564 9940
rect 25620 9884 26348 9940
rect 26404 9884 26414 9940
rect 32834 9884 32844 9940
rect 32900 9884 33852 9940
rect 33908 9884 33918 9940
rect 20514 9772 20524 9828
rect 20580 9772 22204 9828
rect 22260 9772 22270 9828
rect 18162 9660 18172 9716
rect 18228 9660 19068 9716
rect 19124 9660 21308 9716
rect 21364 9660 21374 9716
rect 22764 9604 22820 9884
rect 25890 9772 25900 9828
rect 25956 9772 31388 9828
rect 31444 9772 31454 9828
rect 34178 9772 34188 9828
rect 34244 9772 34748 9828
rect 34804 9772 35980 9828
rect 36036 9772 36046 9828
rect 24770 9660 24780 9716
rect 24836 9660 32284 9716
rect 32340 9660 32350 9716
rect 33282 9660 33292 9716
rect 33348 9660 34524 9716
rect 34580 9660 34590 9716
rect 19170 9548 19180 9604
rect 19236 9548 20076 9604
rect 20132 9548 21252 9604
rect 22754 9548 22764 9604
rect 22820 9548 22830 9604
rect 24434 9548 24444 9604
rect 24500 9548 25228 9604
rect 25284 9548 25294 9604
rect 29586 9548 29596 9604
rect 29652 9548 30380 9604
rect 30436 9548 30446 9604
rect 31938 9548 31948 9604
rect 32004 9548 32396 9604
rect 32452 9548 33068 9604
rect 33124 9548 33134 9604
rect 21196 9492 21252 9548
rect 21196 9436 24332 9492
rect 24388 9436 24398 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 22194 9324 22204 9380
rect 22260 9324 22876 9380
rect 22932 9324 22942 9380
rect 26226 9324 26236 9380
rect 26292 9324 27132 9380
rect 27188 9324 27198 9380
rect 22530 9212 22540 9268
rect 22596 9212 23772 9268
rect 23828 9212 24668 9268
rect 24724 9212 24734 9268
rect 25666 9212 25676 9268
rect 25732 9212 26908 9268
rect 26964 9212 28140 9268
rect 28196 9212 28206 9268
rect 29138 9212 29148 9268
rect 29204 9212 30940 9268
rect 30996 9212 31006 9268
rect 29148 9156 29204 9212
rect 18918 9100 18956 9156
rect 19012 9100 19022 9156
rect 23874 9100 23884 9156
rect 23940 9100 25452 9156
rect 25508 9100 25518 9156
rect 27682 9100 27692 9156
rect 27748 9100 29204 9156
rect 24658 8988 24668 9044
rect 24724 8988 26348 9044
rect 26404 8988 26414 9044
rect 32498 8988 32508 9044
rect 32564 8988 35868 9044
rect 35924 8988 36428 9044
rect 36484 8988 36494 9044
rect 9426 8652 9436 8708
rect 9492 8652 14364 8708
rect 14420 8652 14430 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 15362 8428 15372 8484
rect 15428 8428 16380 8484
rect 16436 8428 18844 8484
rect 18900 8428 19852 8484
rect 19908 8428 19918 8484
rect 28242 8428 28252 8484
rect 28308 8428 29596 8484
rect 29652 8428 29662 8484
rect 6290 8316 6300 8372
rect 6356 8316 8092 8372
rect 8148 8316 10892 8372
rect 10948 8316 11452 8372
rect 11508 8316 13132 8372
rect 13188 8316 13916 8372
rect 13972 8316 13982 8372
rect 19058 8316 19068 8372
rect 19124 8316 20300 8372
rect 20356 8316 20366 8372
rect 20514 8204 20524 8260
rect 20580 8204 21308 8260
rect 21364 8204 22092 8260
rect 22148 8204 22158 8260
rect 41101 8148 41901 8176
rect 14018 8092 14028 8148
rect 14084 8092 14700 8148
rect 14756 8092 14766 8148
rect 16034 8092 16044 8148
rect 16100 8092 19292 8148
rect 19348 8092 21532 8148
rect 21588 8092 21598 8148
rect 22754 8092 22764 8148
rect 22820 8092 24220 8148
rect 24276 8092 24286 8148
rect 40114 8092 40124 8148
rect 40180 8092 41901 8148
rect 22764 8036 22820 8092
rect 41101 8064 41901 8092
rect 19394 7980 19404 8036
rect 19460 7980 21420 8036
rect 21476 7980 22820 8036
rect 26338 7980 26348 8036
rect 26404 7980 27580 8036
rect 27636 7980 28364 8036
rect 28420 7980 28430 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 14354 7756 14364 7812
rect 14420 7756 15036 7812
rect 15092 7756 19684 7812
rect 21634 7756 21644 7812
rect 21700 7756 21980 7812
rect 22036 7756 22428 7812
rect 22484 7756 22494 7812
rect 19628 7700 19684 7756
rect 14914 7644 14924 7700
rect 14980 7644 16044 7700
rect 16100 7644 16110 7700
rect 19628 7644 25452 7700
rect 25508 7644 25518 7700
rect 41101 7476 41901 7504
rect 13122 7420 13132 7476
rect 13188 7420 16492 7476
rect 16548 7420 16558 7476
rect 40002 7420 40012 7476
rect 40068 7420 41901 7476
rect 41101 7392 41901 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 27458 6860 27468 6916
rect 27524 6860 28364 6916
rect 28420 6860 29372 6916
rect 29428 6860 29438 6916
rect 41101 6804 41901 6832
rect 25442 6748 25452 6804
rect 25508 6748 26460 6804
rect 26516 6748 26526 6804
rect 39666 6748 39676 6804
rect 39732 6748 41901 6804
rect 41101 6720 41901 6748
rect 21522 6636 21532 6692
rect 21588 6636 21980 6692
rect 22036 6636 22540 6692
rect 22596 6636 22606 6692
rect 13346 6524 13356 6580
rect 13412 6524 21868 6580
rect 21924 6524 22988 6580
rect 23044 6524 24332 6580
rect 24388 6524 24892 6580
rect 24948 6524 24958 6580
rect 1698 6412 1708 6468
rect 1764 6412 1774 6468
rect 24098 6412 24108 6468
rect 24164 6412 27132 6468
rect 27188 6412 27198 6468
rect 1708 6244 1764 6412
rect 25890 6300 25900 6356
rect 25956 6300 26348 6356
rect 26404 6300 26414 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 924 6188 1764 6244
rect 0 6132 800 6160
rect 924 6132 980 6188
rect 41101 6132 41901 6160
rect 0 6076 980 6132
rect 23202 6076 23212 6132
rect 23268 6076 26012 6132
rect 26068 6076 26078 6132
rect 40114 6076 40124 6132
rect 40180 6076 41901 6132
rect 0 6048 800 6076
rect 41101 6048 41901 6076
rect 23426 5964 23436 6020
rect 23492 5964 24220 6020
rect 24276 5964 24286 6020
rect 38434 5964 38444 6020
rect 38500 5964 39788 6020
rect 39844 5964 39854 6020
rect 25554 5852 25564 5908
rect 25620 5852 28812 5908
rect 28868 5852 32508 5908
rect 32564 5852 32574 5908
rect 39554 5852 39564 5908
rect 39620 5852 40124 5908
rect 40180 5852 40190 5908
rect 0 5460 800 5488
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 41101 5460 41901 5488
rect 0 5404 1708 5460
rect 1764 5404 1774 5460
rect 40114 5404 40124 5460
rect 40180 5404 41901 5460
rect 0 5376 800 5404
rect 41101 5376 41901 5404
rect 21634 5292 21644 5348
rect 21700 5292 23100 5348
rect 23156 5292 26124 5348
rect 26180 5292 26190 5348
rect 25778 5180 25788 5236
rect 25844 5180 26348 5236
rect 26404 5180 26414 5236
rect 18834 5068 18844 5124
rect 18900 5068 19516 5124
rect 19572 5068 22876 5124
rect 22932 5068 22942 5124
rect 24098 5068 24108 5124
rect 24164 5068 26236 5124
rect 26292 5068 26302 5124
rect 1698 4844 1708 4900
rect 1764 4844 1774 4900
rect 0 4788 800 4816
rect 1708 4788 1764 4844
rect 41101 4788 41901 4816
rect 0 4732 1764 4788
rect 40114 4732 40124 4788
rect 40180 4732 41901 4788
rect 0 4704 800 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 41101 4704 41901 4732
rect 19618 4508 19628 4564
rect 19684 4508 19852 4564
rect 19908 4508 19918 4564
rect 0 4116 800 4144
rect 41101 4116 41901 4144
rect 0 4060 1708 4116
rect 1764 4060 1774 4116
rect 40114 4060 40124 4116
rect 40180 4060 41901 4116
rect 0 4032 800 4060
rect 41101 4032 41901 4060
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19506 3612 19516 3668
rect 19572 3612 21196 3668
rect 21252 3612 21262 3668
rect 19282 3500 19292 3556
rect 19348 3500 20748 3556
rect 20804 3500 20814 3556
rect 0 3444 800 3472
rect 41101 3444 41901 3472
rect 0 3388 1708 3444
rect 1764 3388 1774 3444
rect 19618 3388 19628 3444
rect 19684 3388 20188 3444
rect 20244 3388 20254 3444
rect 40124 3388 41901 3444
rect 0 3360 800 3388
rect 40124 3332 40180 3388
rect 41101 3360 41901 3388
rect 40114 3276 40124 3332
rect 40180 3276 40190 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 41101 2772 41901 2800
rect 39666 2716 39676 2772
rect 39732 2716 41901 2772
rect 41101 2688 41901 2716
rect 41101 2100 41901 2128
rect 39218 2044 39228 2100
rect 39284 2044 41901 2100
rect 41101 2016 41901 2044
<< via3 >>
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 17500 35308 17556 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 31164 35084 31220 35140
rect 30156 34524 30212 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 30156 32956 30212 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 18956 31836 19012 31892
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 18956 30940 19012 30996
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 17500 28028 17556 28084
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 31164 25564 31220 25620
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 15484 23212 15540 23268
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 4844 22204 4900 22260
rect 6300 22092 6356 22148
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 7532 21644 7588 21700
rect 33852 21532 33908 21588
rect 15484 21308 15540 21364
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 6300 20524 6356 20580
rect 8540 20524 8596 20580
rect 34524 20524 34580 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 9324 19964 9380 20020
rect 8428 19852 8484 19908
rect 9436 19852 9492 19908
rect 33852 19740 33908 19796
rect 34524 19740 34580 19796
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 4844 19292 4900 19348
rect 8428 19068 8484 19124
rect 19628 19068 19684 19124
rect 31276 19068 31332 19124
rect 17836 18956 17892 19012
rect 19180 18956 19236 19012
rect 18956 18844 19012 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 6300 18508 6356 18564
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 17836 17836 17892 17892
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 7532 16828 7588 16884
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 6300 16156 6356 16212
rect 8540 16156 8596 16212
rect 19292 15820 19348 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 8428 15372 8484 15428
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 9436 14700 9492 14756
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 9324 13692 9380 13748
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 31276 13020 31332 13076
rect 19180 12572 19236 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 18956 9100 19012 9156
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 19628 4508 19684 4564
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19292 3500 19348 3556
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 41580 4768 42396
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 19808 42364 20128 42396
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 17500 35364 17556 35374
rect 17500 28084 17556 35308
rect 19808 34524 20128 36036
rect 35168 41580 35488 42396
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 31164 35140 31220 35150
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 30156 34580 30212 34590
rect 30156 33012 30212 34524
rect 30156 32946 30212 32956
rect 17500 28018 17556 28028
rect 18956 31892 19012 31902
rect 18956 30996 19012 31836
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 15484 23268 15540 23278
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4844 22260 4900 22270
rect 4844 19348 4900 22204
rect 4844 19282 4900 19292
rect 6300 22148 6356 22158
rect 6300 20580 6356 22092
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 6300 18564 6356 20524
rect 6300 16212 6356 18508
rect 7532 21700 7588 21710
rect 7532 16884 7588 21644
rect 15484 21364 15540 23212
rect 15484 21298 15540 21308
rect 8540 20580 8596 20590
rect 7532 16818 7588 16828
rect 8428 19908 8484 19918
rect 8428 19124 8484 19852
rect 6300 16146 6356 16156
rect 8428 15428 8484 19068
rect 8540 16212 8596 20524
rect 8540 16146 8596 16156
rect 9324 20020 9380 20030
rect 8428 15362 8484 15372
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 9324 13748 9380 19964
rect 9436 19908 9492 19918
rect 9436 14756 9492 19852
rect 17836 19012 17892 19022
rect 17836 17892 17892 18956
rect 17836 17826 17892 17836
rect 18956 18900 19012 30940
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 31164 25620 31220 35084
rect 31164 25554 31220 25564
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19628 19124 19684 19134
rect 9436 14690 9492 14700
rect 9324 13682 9380 13692
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 18956 9156 19012 18844
rect 19180 19012 19236 19022
rect 19180 12628 19236 18956
rect 19180 12562 19236 12572
rect 19292 15876 19348 15886
rect 18956 9090 19012 9100
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19292 3556 19348 15820
rect 19628 4564 19684 19068
rect 19628 4498 19684 4508
rect 19808 18844 20128 20356
rect 33852 21588 33908 21598
rect 33852 19796 33908 21532
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 33852 19730 33908 19740
rect 34524 20580 34580 20590
rect 34524 19796 34580 20524
rect 34524 19730 34580 19740
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 31276 19124 31332 19134
rect 31276 13076 31332 19068
rect 31276 13010 31332 13020
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19292 3490 19348 3500
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0553_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0554_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24752 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0555_
timestamp 1698431365
transform -1 0 24080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0556_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22960 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0557_
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0558_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0559_
timestamp 1698431365
transform 1 0 15904 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0560_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0561_
timestamp 1698431365
transform -1 0 16016 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0562_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0563_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0564_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0565_
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0566_
timestamp 1698431365
transform -1 0 38416 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0567_
timestamp 1698431365
transform -1 0 36848 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0568_
timestamp 1698431365
transform 1 0 35056 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0569_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34832 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0570_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26768 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0571_
timestamp 1698431365
transform -1 0 34832 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0572_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0573_
timestamp 1698431365
transform 1 0 12768 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0574_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0575_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0576_
timestamp 1698431365
transform 1 0 17808 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0577_
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0578_
timestamp 1698431365
transform -1 0 24864 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0579_
timestamp 1698431365
transform -1 0 23632 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0580_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22960 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0581_
timestamp 1698431365
transform -1 0 20272 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0582_
timestamp 1698431365
transform -1 0 19488 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0583_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0584_
timestamp 1698431365
transform 1 0 14448 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0585_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0586_
timestamp 1698431365
transform 1 0 18816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0587_
timestamp 1698431365
transform -1 0 19936 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0588_
timestamp 1698431365
transform -1 0 20272 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0589_
timestamp 1698431365
transform -1 0 19488 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0590_
timestamp 1698431365
transform -1 0 16352 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0591_
timestamp 1698431365
transform -1 0 14224 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0592_
timestamp 1698431365
transform -1 0 21840 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0593_
timestamp 1698431365
transform -1 0 17024 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0594_
timestamp 1698431365
transform -1 0 18368 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0595_
timestamp 1698431365
transform -1 0 32144 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0596_
timestamp 1698431365
transform 1 0 30016 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0597_
timestamp 1698431365
transform 1 0 30240 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0598_
timestamp 1698431365
transform -1 0 32704 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0599_
timestamp 1698431365
transform 1 0 29792 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0600_
timestamp 1698431365
transform 1 0 31472 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0601_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31808 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0602_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32032 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0603_
timestamp 1698431365
transform -1 0 30576 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0604_
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0605_
timestamp 1698431365
transform 1 0 32480 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0606_
timestamp 1698431365
transform -1 0 32032 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0607_
timestamp 1698431365
transform -1 0 33936 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0608_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32032 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0609_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0610_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0611_
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0612_
timestamp 1698431365
transform -1 0 30464 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0613_
timestamp 1698431365
transform 1 0 27440 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0614_
timestamp 1698431365
transform -1 0 27776 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0615_
timestamp 1698431365
transform 1 0 17584 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0616_
timestamp 1698431365
transform 1 0 18816 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0617_
timestamp 1698431365
transform -1 0 34272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0618_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0619_
timestamp 1698431365
transform 1 0 34160 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0620_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34496 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0621_
timestamp 1698431365
transform -1 0 34496 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0622_
timestamp 1698431365
transform -1 0 27664 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0623_
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0624_
timestamp 1698431365
transform 1 0 23632 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0625_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0626_
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0627_
timestamp 1698431365
transform -1 0 23968 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0628_
timestamp 1698431365
transform -1 0 26208 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0629_
timestamp 1698431365
transform -1 0 24864 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0630_
timestamp 1698431365
transform -1 0 26544 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0631_
timestamp 1698431365
transform 1 0 25200 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0632_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24192 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0633_
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0634_
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0635_
timestamp 1698431365
transform -1 0 24192 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0636_
timestamp 1698431365
transform 1 0 28448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0637_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0638_
timestamp 1698431365
transform -1 0 28112 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0639_
timestamp 1698431365
transform -1 0 32592 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0640_
timestamp 1698431365
transform -1 0 25536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0641_
timestamp 1698431365
transform 1 0 22288 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0642_
timestamp 1698431365
transform 1 0 24080 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0643_
timestamp 1698431365
transform -1 0 25984 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0644_
timestamp 1698431365
transform 1 0 28112 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0645_
timestamp 1698431365
transform 1 0 28000 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0646_
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0647_
timestamp 1698431365
transform 1 0 29680 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0648_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30352 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0649_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0650_
timestamp 1698431365
transform -1 0 28224 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0651_
timestamp 1698431365
transform -1 0 28448 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0652_
timestamp 1698431365
transform 1 0 26656 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0653_
timestamp 1698431365
transform 1 0 25872 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0654_
timestamp 1698431365
transform -1 0 29680 0 -1 10976
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0655_
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0656_
timestamp 1698431365
transform -1 0 19264 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0657_
timestamp 1698431365
transform 1 0 23968 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0658_
timestamp 1698431365
transform 1 0 23184 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0659_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0660_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0661_
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0662_
timestamp 1698431365
transform 1 0 29008 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0663_
timestamp 1698431365
transform 1 0 17808 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0664_
timestamp 1698431365
transform 1 0 17696 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0665_
timestamp 1698431365
transform 1 0 13328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0666_
timestamp 1698431365
transform 1 0 20384 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0667_
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0668_
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0669_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0670_
timestamp 1698431365
transform -1 0 28448 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0671_
timestamp 1698431365
transform 1 0 31696 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0672_
timestamp 1698431365
transform -1 0 33040 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0673_
timestamp 1698431365
transform -1 0 32592 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0674_
timestamp 1698431365
transform -1 0 34160 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0675_
timestamp 1698431365
transform -1 0 31136 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0676_
timestamp 1698431365
transform -1 0 32592 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0677_
timestamp 1698431365
transform -1 0 37520 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0678_
timestamp 1698431365
transform -1 0 38752 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0679_
timestamp 1698431365
transform -1 0 34832 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0680_
timestamp 1698431365
transform -1 0 31024 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0681_
timestamp 1698431365
transform 1 0 14672 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0682_
timestamp 1698431365
transform 1 0 15680 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0683_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19936 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0684_
timestamp 1698431365
transform -1 0 23968 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0685_
timestamp 1698431365
transform -1 0 21728 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0686_
timestamp 1698431365
transform -1 0 16912 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0687_
timestamp 1698431365
transform 1 0 19488 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0688_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0689_
timestamp 1698431365
transform 1 0 23072 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0690_
timestamp 1698431365
transform -1 0 25984 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0691_
timestamp 1698431365
transform 1 0 30688 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0692_
timestamp 1698431365
transform -1 0 32928 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0693_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34160 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0694_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0695_
timestamp 1698431365
transform -1 0 19824 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0696_
timestamp 1698431365
transform -1 0 20608 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0697_
timestamp 1698431365
transform -1 0 20160 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0698_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0699_
timestamp 1698431365
transform -1 0 20272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0700_
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0701_
timestamp 1698431365
transform 1 0 9632 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0702_
timestamp 1698431365
transform -1 0 15456 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0703_
timestamp 1698431365
transform -1 0 14784 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0704_
timestamp 1698431365
transform -1 0 21504 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0705_
timestamp 1698431365
transform 1 0 19824 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0706_
timestamp 1698431365
transform 1 0 21728 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0707_
timestamp 1698431365
transform 1 0 23632 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0708_
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0709_
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0710_
timestamp 1698431365
transform -1 0 20720 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0711_
timestamp 1698431365
transform 1 0 21840 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0712_
timestamp 1698431365
transform 1 0 24528 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0713_
timestamp 1698431365
transform -1 0 27104 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0714_
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0715_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0716_
timestamp 1698431365
transform 1 0 25984 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0717_
timestamp 1698431365
transform 1 0 22960 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0718_
timestamp 1698431365
transform 1 0 24080 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0719_
timestamp 1698431365
transform -1 0 24528 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0720_
timestamp 1698431365
transform 1 0 23520 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0721_
timestamp 1698431365
transform 1 0 25088 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0722_
timestamp 1698431365
transform -1 0 10640 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0723_
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0724_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0725_
timestamp 1698431365
transform 1 0 3472 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0726_
timestamp 1698431365
transform -1 0 3360 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0727_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3808 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0728_
timestamp 1698431365
transform 1 0 8512 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0729_
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0730_
timestamp 1698431365
transform 1 0 11984 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0731_
timestamp 1698431365
transform -1 0 12320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0732_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0733_
timestamp 1698431365
transform -1 0 10976 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0734_
timestamp 1698431365
transform 1 0 8288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0735_
timestamp 1698431365
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0736_
timestamp 1698431365
transform 1 0 9520 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0737_
timestamp 1698431365
transform 1 0 8288 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0738_
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0739_
timestamp 1698431365
transform 1 0 6496 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0740_
timestamp 1698431365
transform 1 0 3584 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0741_
timestamp 1698431365
transform 1 0 2800 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0742_
timestamp 1698431365
transform 1 0 4032 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0743_
timestamp 1698431365
transform 1 0 6384 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0744_
timestamp 1698431365
transform 1 0 7056 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0745_
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0746_
timestamp 1698431365
transform -1 0 7840 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0747_
timestamp 1698431365
transform 1 0 7840 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0748_
timestamp 1698431365
transform 1 0 11088 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0749_
timestamp 1698431365
transform 1 0 9408 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0750_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0751_
timestamp 1698431365
transform 1 0 6160 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0752_
timestamp 1698431365
transform 1 0 10752 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0753_
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0754_
timestamp 1698431365
transform -1 0 8288 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0755_
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0756_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0757_
timestamp 1698431365
transform 1 0 7728 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0758_
timestamp 1698431365
transform 1 0 3360 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0759_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0760_
timestamp 1698431365
transform 1 0 5936 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0761_
timestamp 1698431365
transform 1 0 9408 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0762_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7280 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0763_
timestamp 1698431365
transform -1 0 24416 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0764_
timestamp 1698431365
transform -1 0 9408 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0765_
timestamp 1698431365
transform -1 0 8624 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0766_
timestamp 1698431365
transform -1 0 10528 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0767_
timestamp 1698431365
transform -1 0 7280 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0768_
timestamp 1698431365
transform 1 0 5376 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0769_
timestamp 1698431365
transform 1 0 5600 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0770_
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0771_
timestamp 1698431365
transform -1 0 8848 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0772_
timestamp 1698431365
transform 1 0 8512 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0773_
timestamp 1698431365
transform -1 0 23072 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0774_
timestamp 1698431365
transform -1 0 6720 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0775_
timestamp 1698431365
transform 1 0 4256 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0776_
timestamp 1698431365
transform 1 0 11424 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0777_
timestamp 1698431365
transform -1 0 6608 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0778_
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0779_
timestamp 1698431365
transform -1 0 8064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0780_
timestamp 1698431365
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0781_
timestamp 1698431365
transform -1 0 5264 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0782_
timestamp 1698431365
transform 1 0 5488 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0783_
timestamp 1698431365
transform 1 0 6048 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0784_
timestamp 1698431365
transform 1 0 6608 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0785_
timestamp 1698431365
transform 1 0 6944 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0786_
timestamp 1698431365
transform -1 0 8288 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0787_
timestamp 1698431365
transform -1 0 3808 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0788_
timestamp 1698431365
transform -1 0 26880 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0789_
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0790_
timestamp 1698431365
transform -1 0 10416 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0791_
timestamp 1698431365
transform 1 0 2912 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0792_
timestamp 1698431365
transform 1 0 6160 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0793_
timestamp 1698431365
transform 1 0 7056 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0794_
timestamp 1698431365
transform -1 0 8064 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0795_
timestamp 1698431365
transform 1 0 5936 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0796_
timestamp 1698431365
transform 1 0 6720 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0797_
timestamp 1698431365
transform 1 0 7840 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0798_
timestamp 1698431365
transform 1 0 8064 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0799_
timestamp 1698431365
transform -1 0 9856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0800_
timestamp 1698431365
transform 1 0 10528 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0801_
timestamp 1698431365
transform 1 0 4368 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0802_
timestamp 1698431365
transform -1 0 7168 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0803_
timestamp 1698431365
transform -1 0 5936 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0804_
timestamp 1698431365
transform -1 0 5264 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0805_
timestamp 1698431365
transform -1 0 7056 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0806_
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0807_
timestamp 1698431365
transform 1 0 4592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0808_
timestamp 1698431365
transform -1 0 6944 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0809_
timestamp 1698431365
transform 1 0 4816 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0810_
timestamp 1698431365
transform 1 0 21728 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0811_
timestamp 1698431365
transform -1 0 8176 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0812_
timestamp 1698431365
transform 1 0 7056 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0813_
timestamp 1698431365
transform -1 0 4368 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0814_
timestamp 1698431365
transform 1 0 4816 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0815_
timestamp 1698431365
transform -1 0 6496 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0816_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0817_
timestamp 1698431365
transform 1 0 5488 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0818_
timestamp 1698431365
transform 1 0 5376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0819_
timestamp 1698431365
transform 1 0 4256 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0820_
timestamp 1698431365
transform -1 0 6944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0821_
timestamp 1698431365
transform 1 0 5040 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0822_
timestamp 1698431365
transform 1 0 6272 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0823_
timestamp 1698431365
transform -1 0 7056 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0824_
timestamp 1698431365
transform -1 0 4368 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0825_
timestamp 1698431365
transform -1 0 12880 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0826_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0827_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0828_
timestamp 1698431365
transform -1 0 10304 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0829_
timestamp 1698431365
transform 1 0 22400 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0830_
timestamp 1698431365
transform 1 0 23968 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0831_
timestamp 1698431365
transform -1 0 10752 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0832_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0833_
timestamp 1698431365
transform 1 0 7728 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0834_
timestamp 1698431365
transform -1 0 6160 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0835_
timestamp 1698431365
transform 1 0 7952 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0836_
timestamp 1698431365
transform 1 0 8512 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0837_
timestamp 1698431365
transform 1 0 11200 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0838_
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0839_
timestamp 1698431365
transform -1 0 10304 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0840_
timestamp 1698431365
transform 1 0 9184 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0841_
timestamp 1698431365
transform -1 0 10080 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0842_
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0843_
timestamp 1698431365
transform -1 0 8288 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0844_
timestamp 1698431365
transform 1 0 10640 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0845_
timestamp 1698431365
transform -1 0 22624 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0846_
timestamp 1698431365
transform 1 0 12544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0847_
timestamp 1698431365
transform 1 0 13104 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0848_
timestamp 1698431365
transform 1 0 9968 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0849_
timestamp 1698431365
transform -1 0 11872 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0850_
timestamp 1698431365
transform 1 0 9520 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0851_
timestamp 1698431365
transform -1 0 12208 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0852_
timestamp 1698431365
transform -1 0 23856 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0853_
timestamp 1698431365
transform -1 0 12880 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0854_
timestamp 1698431365
transform -1 0 10080 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0855_
timestamp 1698431365
transform 1 0 11536 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0856_
timestamp 1698431365
transform -1 0 11312 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0857_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12544 0 -1 34496
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0858_
timestamp 1698431365
transform -1 0 14672 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0859_
timestamp 1698431365
transform 1 0 12880 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0860_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0861_
timestamp 1698431365
transform -1 0 12880 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0862_
timestamp 1698431365
transform 1 0 15456 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0863_
timestamp 1698431365
transform 1 0 15344 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0864_
timestamp 1698431365
transform -1 0 16016 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0865_
timestamp 1698431365
transform -1 0 16912 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0866_
timestamp 1698431365
transform -1 0 18032 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0867_
timestamp 1698431365
transform -1 0 16800 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0868_
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0869_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0870_
timestamp 1698431365
transform -1 0 16576 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0871_
timestamp 1698431365
transform -1 0 15344 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0872_
timestamp 1698431365
transform 1 0 14560 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0873_
timestamp 1698431365
transform 1 0 15008 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0874_
timestamp 1698431365
transform -1 0 15232 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0875_
timestamp 1698431365
transform 1 0 15904 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0876_
timestamp 1698431365
transform -1 0 14000 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0877_
timestamp 1698431365
transform 1 0 22736 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0878_
timestamp 1698431365
transform 1 0 18704 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0879_
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0880_
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0881_
timestamp 1698431365
transform -1 0 22176 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0882_
timestamp 1698431365
transform -1 0 21840 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0883_
timestamp 1698431365
transform -1 0 26992 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0884_
timestamp 1698431365
transform -1 0 24528 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0885_
timestamp 1698431365
transform 1 0 23632 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0886_
timestamp 1698431365
transform -1 0 26320 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0887_
timestamp 1698431365
transform -1 0 29680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0888_
timestamp 1698431365
transform 1 0 25536 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0889_
timestamp 1698431365
transform -1 0 26096 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0890_
timestamp 1698431365
transform 1 0 24528 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0891_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0892_
timestamp 1698431365
transform -1 0 29680 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0893_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0894_
timestamp 1698431365
transform 1 0 26320 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0895_
timestamp 1698431365
transform -1 0 27776 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0896_
timestamp 1698431365
transform 1 0 27664 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0897_
timestamp 1698431365
transform 1 0 24864 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0898_
timestamp 1698431365
transform -1 0 28784 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0899_
timestamp 1698431365
transform -1 0 27776 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0900_
timestamp 1698431365
transform 1 0 30352 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0901_
timestamp 1698431365
transform 1 0 32032 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1698431365
transform 1 0 31584 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0903_
timestamp 1698431365
transform 1 0 30128 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0904_
timestamp 1698431365
transform 1 0 29792 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _0905_
timestamp 1698431365
transform -1 0 31920 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0906_
timestamp 1698431365
transform -1 0 31696 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0907_
timestamp 1698431365
transform 1 0 31696 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0908_
timestamp 1698431365
transform 1 0 30016 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0909_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0910_
timestamp 1698431365
transform -1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0911_
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0912_
timestamp 1698431365
transform 1 0 29232 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0913_
timestamp 1698431365
transform -1 0 34272 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0914_
timestamp 1698431365
transform -1 0 33376 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0915_
timestamp 1698431365
transform -1 0 32704 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0916_
timestamp 1698431365
transform -1 0 31696 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0917_
timestamp 1698431365
transform 1 0 30688 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0918_
timestamp 1698431365
transform -1 0 31584 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _0919_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31024 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0920_
timestamp 1698431365
transform -1 0 32480 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0921_
timestamp 1698431365
transform -1 0 30688 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0922_
timestamp 1698431365
transform 1 0 31024 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0923_
timestamp 1698431365
transform 1 0 28784 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0924_
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0925_
timestamp 1698431365
transform 1 0 24192 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0926_
timestamp 1698431365
transform 1 0 25424 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0927_
timestamp 1698431365
transform 1 0 22624 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0928_
timestamp 1698431365
transform -1 0 36512 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0929_
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0930_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30576 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0931_
timestamp 1698431365
transform 1 0 36064 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0932_
timestamp 1698431365
transform -1 0 36064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0933_
timestamp 1698431365
transform -1 0 37968 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0934_
timestamp 1698431365
transform -1 0 37520 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0935_
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0936_
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0937_
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0938_
timestamp 1698431365
transform -1 0 36848 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0939_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0940_
timestamp 1698431365
transform -1 0 35168 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0941_
timestamp 1698431365
transform -1 0 36512 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0942_
timestamp 1698431365
transform 1 0 35168 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0943_
timestamp 1698431365
transform 1 0 37520 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0944_
timestamp 1698431365
transform -1 0 27216 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0945_
timestamp 1698431365
transform -1 0 34944 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0946_
timestamp 1698431365
transform -1 0 33600 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0947_
timestamp 1698431365
transform 1 0 29680 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0948_
timestamp 1698431365
transform -1 0 28672 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0949_
timestamp 1698431365
transform 1 0 26432 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0950_
timestamp 1698431365
transform -1 0 28224 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0951_
timestamp 1698431365
transform -1 0 26880 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0952_
timestamp 1698431365
transform 1 0 25760 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0953_
timestamp 1698431365
transform 1 0 22624 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0954_
timestamp 1698431365
transform -1 0 29792 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0955_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0956_
timestamp 1698431365
transform 1 0 11648 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0957_
timestamp 1698431365
transform -1 0 14448 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0958_
timestamp 1698431365
transform -1 0 14672 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0959_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0960_
timestamp 1698431365
transform -1 0 14672 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _0961_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13552 0 -1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0962_
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0963_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16128 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0964_
timestamp 1698431365
transform -1 0 15904 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0965_
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0966_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0967_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0968_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0969_
timestamp 1698431365
transform 1 0 13440 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0970_
timestamp 1698431365
transform 1 0 11872 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0971_
timestamp 1698431365
transform 1 0 12768 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0972_
timestamp 1698431365
transform 1 0 13552 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0973_
timestamp 1698431365
transform 1 0 14672 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0974_
timestamp 1698431365
transform -1 0 24640 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0975_
timestamp 1698431365
transform 1 0 31808 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0976_
timestamp 1698431365
transform 1 0 30464 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0977_
timestamp 1698431365
transform -1 0 33152 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0978_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0979_
timestamp 1698431365
transform -1 0 37520 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0980_
timestamp 1698431365
transform -1 0 34496 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0981_
timestamp 1698431365
transform -1 0 33824 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0982_
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0983_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0984_
timestamp 1698431365
transform -1 0 32480 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0985_
timestamp 1698431365
transform 1 0 35280 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0986_
timestamp 1698431365
transform -1 0 39200 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0987_
timestamp 1698431365
transform -1 0 36624 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0988_
timestamp 1698431365
transform 1 0 26880 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0989_
timestamp 1698431365
transform 1 0 25536 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0990_
timestamp 1698431365
transform 1 0 27104 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0991_
timestamp 1698431365
transform -1 0 33488 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0992_
timestamp 1698431365
transform 1 0 35504 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0993_
timestamp 1698431365
transform -1 0 36176 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0994_
timestamp 1698431365
transform -1 0 36512 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0995_
timestamp 1698431365
transform -1 0 33712 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0996_
timestamp 1698431365
transform 1 0 31248 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0997_
timestamp 1698431365
transform -1 0 35952 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0998_
timestamp 1698431365
transform -1 0 35056 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0999_
timestamp 1698431365
transform -1 0 32592 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1000_
timestamp 1698431365
transform 1 0 31696 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1001_
timestamp 1698431365
transform 1 0 28224 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1002_
timestamp 1698431365
transform 1 0 29344 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1003_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1004_
timestamp 1698431365
transform -1 0 19488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1005_
timestamp 1698431365
transform -1 0 18816 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1006_
timestamp 1698431365
transform 1 0 17024 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1007_
timestamp 1698431365
transform -1 0 14448 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1008_
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1009_
timestamp 1698431365
transform 1 0 29680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1010_
timestamp 1698431365
transform -1 0 27888 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1011_
timestamp 1698431365
transform 1 0 18704 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1012_
timestamp 1698431365
transform 1 0 16464 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1013_
timestamp 1698431365
transform 1 0 14448 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1014_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1015_
timestamp 1698431365
transform 1 0 11760 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1016_
timestamp 1698431365
transform 1 0 10864 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1017_
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1018_
timestamp 1698431365
transform -1 0 21616 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1019_
timestamp 1698431365
transform 1 0 15344 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1020_
timestamp 1698431365
transform 1 0 15680 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1021_
timestamp 1698431365
transform -1 0 19264 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1022_
timestamp 1698431365
transform 1 0 17584 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1023_
timestamp 1698431365
transform 1 0 19264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1024_
timestamp 1698431365
transform -1 0 19936 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1025_
timestamp 1698431365
transform 1 0 18256 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1026_
timestamp 1698431365
transform -1 0 20160 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1027_
timestamp 1698431365
transform 1 0 19712 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1028_
timestamp 1698431365
transform -1 0 22400 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1029_
timestamp 1698431365
transform 1 0 15680 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1030_
timestamp 1698431365
transform 1 0 18032 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1031_
timestamp 1698431365
transform 1 0 18032 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1032_
timestamp 1698431365
transform 1 0 18480 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1033_
timestamp 1698431365
transform -1 0 19376 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1034_
timestamp 1698431365
transform -1 0 18032 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1035_
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1036_
timestamp 1698431365
transform -1 0 19376 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1037_
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1038_
timestamp 1698431365
transform 1 0 19040 0 -1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1039_
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1040_
timestamp 1698431365
transform 1 0 32816 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1041_
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1042_
timestamp 1698431365
transform -1 0 37632 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1043_
timestamp 1698431365
transform -1 0 34384 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1044_
timestamp 1698431365
transform 1 0 32144 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698431365
transform 1 0 34384 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1046_
timestamp 1698431365
transform -1 0 22624 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1047_
timestamp 1698431365
transform 1 0 31360 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1048_
timestamp 1698431365
transform -1 0 31360 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1049_
timestamp 1698431365
transform 1 0 32480 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1050_
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1051_
timestamp 1698431365
transform -1 0 32704 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1052_
timestamp 1698431365
transform 1 0 33376 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1053_
timestamp 1698431365
transform 1 0 34832 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1054_
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1055_
timestamp 1698431365
transform -1 0 34944 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1056_
timestamp 1698431365
transform 1 0 35168 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1057_
timestamp 1698431365
transform 1 0 36400 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1058_
timestamp 1698431365
transform -1 0 35168 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1059_
timestamp 1698431365
transform 1 0 33600 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1060_
timestamp 1698431365
transform 1 0 35952 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1061_
timestamp 1698431365
transform 1 0 35728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1062_
timestamp 1698431365
transform -1 0 36400 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1063_
timestamp 1698431365
transform 1 0 36848 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1064_
timestamp 1698431365
transform 1 0 36736 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1065_
timestamp 1698431365
transform 1 0 37632 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1066_
timestamp 1698431365
transform -1 0 38752 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1067_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1068_
timestamp 1698431365
transform -1 0 37856 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1069_
timestamp 1698431365
transform 1 0 11200 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1070_
timestamp 1698431365
transform 1 0 9856 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1071_
timestamp 1698431365
transform 1 0 10416 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1072_
timestamp 1698431365
transform -1 0 14784 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1073_
timestamp 1698431365
transform 1 0 11648 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1074_
timestamp 1698431365
transform 1 0 11872 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1075_
timestamp 1698431365
transform 1 0 13552 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1076_
timestamp 1698431365
transform -1 0 25088 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1077_
timestamp 1698431365
transform 1 0 25200 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1078_
timestamp 1698431365
transform 1 0 15456 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1079_
timestamp 1698431365
transform -1 0 18928 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1080_
timestamp 1698431365
transform -1 0 16800 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1081_
timestamp 1698431365
transform -1 0 21840 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1082_
timestamp 1698431365
transform -1 0 18368 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1083_
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1084_
timestamp 1698431365
transform -1 0 20832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1085_
timestamp 1698431365
transform 1 0 16240 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1086_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1087_
timestamp 1698431365
transform 1 0 16688 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1088_
timestamp 1698431365
transform -1 0 18928 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1089_
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1090_
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1091_
timestamp 1698431365
transform -1 0 18480 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1092_
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1093_
timestamp 1698431365
transform 1 0 18928 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1094_
timestamp 1698431365
transform 1 0 19264 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1095_
timestamp 1698431365
transform 1 0 21952 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1096_
timestamp 1698431365
transform -1 0 17024 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1097_
timestamp 1698431365
transform -1 0 18816 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1098_
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1099_
timestamp 1698431365
transform 1 0 16464 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1100_
timestamp 1698431365
transform 1 0 17808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1101_
timestamp 1698431365
transform 1 0 17360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1102_
timestamp 1698431365
transform -1 0 17808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1103_
timestamp 1698431365
transform -1 0 17696 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1104_
timestamp 1698431365
transform 1 0 17360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1105_
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1106_
timestamp 1698431365
transform 1 0 16016 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1107_
timestamp 1698431365
transform -1 0 15904 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1108_
timestamp 1698431365
transform 1 0 17696 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1109_
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1110_
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1111_
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1112_
timestamp 1698431365
transform 1 0 21280 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1113_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1114_
timestamp 1698431365
transform 1 0 18592 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1115_
timestamp 1698431365
transform 1 0 19264 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1116_
timestamp 1698431365
transform 1 0 22736 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1117_
timestamp 1698431365
transform 1 0 25312 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1118_
timestamp 1698431365
transform 1 0 10752 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1119_
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1120_
timestamp 1698431365
transform 1 0 2128 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1121_
timestamp 1698431365
transform 1 0 1792 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1122_
timestamp 1698431365
transform 1 0 7952 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1123_
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1124_
timestamp 1698431365
transform -1 0 11648 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1125_
timestamp 1698431365
transform -1 0 4816 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1126_
timestamp 1698431365
transform -1 0 4816 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1127_
timestamp 1698431365
transform 1 0 6160 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1128_
timestamp 1698431365
transform 1 0 4480 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1129_
timestamp 1698431365
transform -1 0 8736 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1130_
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1131_
timestamp 1698431365
transform 1 0 11088 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1132_
timestamp 1698431365
transform -1 0 19376 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1133_
timestamp 1698431365
transform 1 0 11984 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1134_
timestamp 1698431365
transform -1 0 22736 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1135_
timestamp 1698431365
transform 1 0 22848 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1136_
timestamp 1698431365
transform 1 0 23296 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1137_
timestamp 1698431365
transform 1 0 25648 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1138_
timestamp 1698431365
transform 1 0 29456 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1139_
timestamp 1698431365
transform 1 0 31472 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1140_
timestamp 1698431365
transform 1 0 24864 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1141_
timestamp 1698431365
transform 1 0 37072 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1142_
timestamp 1698431365
transform 1 0 37072 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1143_
timestamp 1698431365
transform 1 0 24976 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1144_
timestamp 1698431365
transform -1 0 26096 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1145_
timestamp 1698431365
transform 1 0 27440 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1146_
timestamp 1698431365
transform -1 0 13888 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1147_
timestamp 1698431365
transform 1 0 26432 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1148_
timestamp 1698431365
transform -1 0 24416 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1149_
timestamp 1698431365
transform -1 0 36624 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1150_
timestamp 1698431365
transform -1 0 36176 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1151_
timestamp 1698431365
transform -1 0 32704 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1152_
timestamp 1698431365
transform -1 0 36624 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1153_
timestamp 1698431365
transform -1 0 36624 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1154_
timestamp 1698431365
transform 1 0 37072 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1155_ asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1156_
timestamp 1698431365
transform 1 0 37072 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1157_
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1158_
timestamp 1698431365
transform 1 0 37072 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1159_
timestamp 1698431365
transform 1 0 25088 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1160_
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1161_
timestamp 1698431365
transform 1 0 19712 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1162_
timestamp 1698431365
transform 1 0 16128 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1163_
timestamp 1698431365
transform 1 0 21616 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1164_
timestamp 1698431365
transform -1 0 16464 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1165_
timestamp 1698431365
transform 1 0 11424 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1166_
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1167_
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1168_
timestamp 1698431365
transform -1 0 23968 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1169_
timestamp 1698431365
transform 1 0 21280 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1202_
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1203_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1204_
timestamp 1698431365
transform 1 0 31696 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1205_
timestamp 1698431365
transform 1 0 29344 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1206_
timestamp 1698431365
transform 1 0 31472 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1207_
timestamp 1698431365
transform 1 0 29680 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1208_
timestamp 1698431365
transform 1 0 30352 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__I asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0585__A1
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0589__A1
timestamp 1698431365
transform -1 0 19936 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0596__I
timestamp 1698431365
transform 1 0 29792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0598__I
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0626__A1
timestamp 1698431365
transform 1 0 22848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0643__A2
timestamp 1698431365
transform -1 0 26208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0649__A1
timestamp 1698431365
transform 1 0 25088 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0652__A2
timestamp 1698431365
transform 1 0 29120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0691__A1
timestamp 1698431365
transform 1 0 31920 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0691__A3
timestamp 1698431365
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0695__I
timestamp 1698431365
transform 1 0 18928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0696__A2
timestamp 1698431365
transform 1 0 21056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A2
timestamp 1698431365
transform -1 0 14112 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0703__A1
timestamp 1698431365
transform 1 0 15008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0705__A2
timestamp 1698431365
transform 1 0 20944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0706__I
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0708__A2
timestamp 1698431365
transform -1 0 18816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0709__A3
timestamp 1698431365
transform -1 0 21168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0710__A1
timestamp 1698431365
transform -1 0 19824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0714__B
timestamp 1698431365
transform 1 0 22960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0718__A1
timestamp 1698431365
transform 1 0 24864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0721__A1
timestamp 1698431365
transform 1 0 26432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0730__A1
timestamp 1698431365
transform -1 0 11984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0730__B
timestamp 1698431365
transform 1 0 13328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0734__A1
timestamp 1698431365
transform -1 0 8288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0734__B
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0736__B
timestamp 1698431365
transform -1 0 10864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__C
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0749__A2
timestamp 1698431365
transform 1 0 10528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0750__A1
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0753__A1
timestamp 1698431365
transform 1 0 9184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0764__B2
timestamp 1698431365
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A1
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0772__A1
timestamp 1698431365
transform 1 0 9408 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__I
timestamp 1698431365
transform 1 0 6944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__B2
timestamp 1698431365
transform 1 0 8512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__B
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0800__A1
timestamp 1698431365
transform 1 0 11424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0810__I
timestamp 1698431365
transform -1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0811__I
timestamp 1698431365
transform -1 0 8400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__A2
timestamp 1698431365
transform 1 0 10528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__B
timestamp 1698431365
transform 1 0 10976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A2
timestamp 1698431365
transform 1 0 10864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698431365
transform 1 0 21504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__A2
timestamp 1698431365
transform 1 0 8960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__I
timestamp 1698431365
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__A2
timestamp 1698431365
transform 1 0 9184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__I
timestamp 1698431365
transform 1 0 22960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A1
timestamp 1698431365
transform 1 0 16800 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A2
timestamp 1698431365
transform 1 0 16352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__A1
timestamp 1698431365
transform 1 0 18032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__B
timestamp 1698431365
transform -1 0 14336 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__I
timestamp 1698431365
transform 1 0 22512 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__A2
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__B
timestamp 1698431365
transform -1 0 24976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__A2
timestamp 1698431365
transform 1 0 23408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A2
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__A2
timestamp 1698431365
transform 1 0 28000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__B2
timestamp 1698431365
transform 1 0 27328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__A2
timestamp 1698431365
transform -1 0 30912 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__B2
timestamp 1698431365
transform -1 0 30464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A2
timestamp 1698431365
transform 1 0 29008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__A1
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__B
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__B
timestamp 1698431365
transform 1 0 31808 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A2
timestamp 1698431365
transform 1 0 23968 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__B
timestamp 1698431365
transform 1 0 27328 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__I
timestamp 1698431365
transform 1 0 22400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__B
timestamp 1698431365
transform 1 0 34944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__A2
timestamp 1698431365
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A1
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__B2
timestamp 1698431365
transform -1 0 35168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__A1
timestamp 1698431365
transform 1 0 38416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__A2
timestamp 1698431365
transform -1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__A1
timestamp 1698431365
transform 1 0 25872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__B
timestamp 1698431365
transform 1 0 26880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__A1
timestamp 1698431365
transform -1 0 21952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0965__A1
timestamp 1698431365
transform 1 0 15344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A1
timestamp 1698431365
transform -1 0 28672 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__A1
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A1
timestamp 1698431365
transform 1 0 14448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__A1
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A1
timestamp 1698431365
transform -1 0 12432 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A1
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A1
timestamp 1698431365
transform 1 0 19376 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A1
timestamp 1698431365
transform 1 0 19936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A1
timestamp 1698431365
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A2
timestamp 1698431365
transform 1 0 30128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A1
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A1
timestamp 1698431365
transform -1 0 33936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698431365
transform 1 0 33152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698431365
transform 1 0 24976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__A1
timestamp 1698431365
transform -1 0 20384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A2
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__I
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A3
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A1
timestamp 1698431365
transform 1 0 17584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A1
timestamp 1698431365
transform -1 0 20832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A1
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__A1
timestamp 1698431365
transform 1 0 17024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__A2
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A1
timestamp 1698431365
transform 1 0 18256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__C
timestamp 1698431365
transform 1 0 17808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__B
timestamp 1698431365
transform 1 0 18928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A1
timestamp 1698431365
transform 1 0 18480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__CLK
timestamp 1698431365
transform 1 0 16464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__CLK
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__CLK
timestamp 1698431365
transform 1 0 14000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__CLK
timestamp 1698431365
transform 1 0 6272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__CLK
timestamp 1698431365
transform 1 0 4480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__CLK
timestamp 1698431365
transform 1 0 11424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__CLK
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1132__CLK
timestamp 1698431365
transform 1 0 19600 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__CLK
timestamp 1698431365
transform 1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__CLK
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__CLK
timestamp 1698431365
transform 1 0 26768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__CLK
timestamp 1698431365
transform -1 0 29456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__CLK
timestamp 1698431365
transform 1 0 31248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__CLK
timestamp 1698431365
transform -1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__CLK
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__CLK
timestamp 1698431365
transform 1 0 36848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__CLK
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__CLK
timestamp 1698431365
transform 1 0 26096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__CLK
timestamp 1698431365
transform 1 0 30912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__CLK
timestamp 1698431365
transform -1 0 29904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__CLK
timestamp 1698431365
transform 1 0 24640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__CLK
timestamp 1698431365
transform 1 0 36848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__CLK
timestamp 1698431365
transform 1 0 32816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__CLK
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__CLK
timestamp 1698431365
transform 1 0 36848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__CLK
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__CLK
timestamp 1698431365
transform 1 0 36176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__CLK
timestamp 1698431365
transform -1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__CLK
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__CLK
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__CLK
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__CLK
timestamp 1698431365
transform 1 0 25536 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__CLK
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1169__CLK
timestamp 1698431365
transform 1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 23184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 18928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 26656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 16800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 26880 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_wb_clk_i_I
timestamp 1698431365
transform -1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout26_I
timestamp 1698431365
transform 1 0 29904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 39648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 39648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 19712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 39648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 23184 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 18928 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1698431365
transform 1 0 27104 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1698431365
transform -1 0 16128 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1698431365
transform -1 0 16800 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1698431365
transform 1 0 27104 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1698431365
transform 1 0 25200 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout22
timestamp 1698431365
transform 1 0 31024 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout23
timestamp 1698431365
transform -1 0 30352 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout24
timestamp 1698431365
transform -1 0 31024 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout25
timestamp 1698431365
transform -1 0 31472 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout26
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout27
timestamp 1698431365
transform 1 0 25424 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_6 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_22 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_30 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_78 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_83 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_89
timestamp 1698431365
transform 1 0 11312 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_97
timestamp 1698431365
transform 1 0 12208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_154
timestamp 1698431365
transform 1 0 18592 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_182
timestamp 1698431365
transform 1 0 21728 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698431365
transform 1 0 23968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_282
timestamp 1698431365
transform 1 0 32928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_287
timestamp 1698431365
transform 1 0 33488 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_324
timestamp 1698431365
transform 1 0 37632 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_332
timestamp 1698431365
transform 1 0 38528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_6 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_158
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_189
timestamp 1698431365
transform 1 0 22512 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_197
timestamp 1698431365
transform 1 0 23408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698431365
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698431365
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698431365
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_330
timestamp 1698431365
transform 1 0 38304 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_338
timestamp 1698431365
transform 1 0 39200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6
timestamp 1698431365
transform 1 0 2016 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698431365
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698431365
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_183
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_242
timestamp 1698431365
transform 1 0 28448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_335
timestamp 1698431365
transform 1 0 38864 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_343
timestamp 1698431365
transform 1 0 39760 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_6
timestamp 1698431365
transform 1 0 2016 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_191
timestamp 1698431365
transform 1 0 22736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_243
timestamp 1698431365
transform 1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_247
timestamp 1698431365
transform 1 0 29008 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_330
timestamp 1698431365
transform 1 0 38304 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_338
timestamp 1698431365
transform 1 0 39200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_6
timestamp 1698431365
transform 1 0 2016 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_22
timestamp 1698431365
transform 1 0 3808 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_30
timestamp 1698431365
transform 1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_195
timestamp 1698431365
transform 1 0 23184 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_208
timestamp 1698431365
transform 1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_222
timestamp 1698431365
transform 1 0 26208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_226
timestamp 1698431365
transform 1 0 26656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_228
timestamp 1698431365
transform 1 0 26880 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_235
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_333
timestamp 1698431365
transform 1 0 38640 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_341
timestamp 1698431365
transform 1 0 39536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_343
timestamp 1698431365
transform 1 0 39760 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_133
timestamp 1698431365
transform 1 0 16240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_137
timestamp 1698431365
transform 1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_174
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_177
timestamp 1698431365
transform 1 0 21168 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_338
timestamp 1698431365
transform 1 0 39200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_53
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_57
timestamp 1698431365
transform 1 0 7728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_88
timestamp 1698431365
transform 1 0 11200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_92
timestamp 1698431365
transform 1 0 11648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_100
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_111
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_120
timestamp 1698431365
transform 1 0 14784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_124
timestamp 1698431365
transform 1 0 15232 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_161
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_173
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_193
timestamp 1698431365
transform 1 0 22960 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_217
timestamp 1698431365
transform 1 0 25648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_219
timestamp 1698431365
transform 1 0 25872 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_222
timestamp 1698431365
transform 1 0 26208 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_230
timestamp 1698431365
transform 1 0 27104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_232
timestamp 1698431365
transform 1 0 27328 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_271
timestamp 1698431365
transform 1 0 31696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_279
timestamp 1698431365
transform 1 0 32592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_283
timestamp 1698431365
transform 1 0 33040 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_333
timestamp 1698431365
transform 1 0 38640 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_80
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_113
timestamp 1698431365
transform 1 0 14000 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_126
timestamp 1698431365
transform 1 0 15456 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_134
timestamp 1698431365
transform 1 0 16352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_193
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_197
timestamp 1698431365
transform 1 0 23408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_203
timestamp 1698431365
transform 1 0 24080 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_225
timestamp 1698431365
transform 1 0 26544 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_246
timestamp 1698431365
transform 1 0 28896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_250
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_311
timestamp 1698431365
transform 1 0 36176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_315
timestamp 1698431365
transform 1 0 36624 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_347
timestamp 1698431365
transform 1 0 40208 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_63
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_70
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_74
timestamp 1698431365
transform 1 0 9632 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_90
timestamp 1698431365
transform 1 0 11424 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_98
timestamp 1698431365
transform 1 0 12320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_115
timestamp 1698431365
transform 1 0 14224 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_160
timestamp 1698431365
transform 1 0 19264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_162
timestamp 1698431365
transform 1 0 19488 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_190
timestamp 1698431365
transform 1 0 22624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_202
timestamp 1698431365
transform 1 0 23968 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_216
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_218
timestamp 1698431365
transform 1 0 25760 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_242
timestamp 1698431365
transform 1 0 28448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_253
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_257
timestamp 1698431365
transform 1 0 30128 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_266
timestamp 1698431365
transform 1 0 31136 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_287
timestamp 1698431365
transform 1 0 33488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_301
timestamp 1698431365
transform 1 0 35056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_333
timestamp 1698431365
transform 1 0 38640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_341
timestamp 1698431365
transform 1 0 39536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_345
timestamp 1698431365
transform 1 0 39984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_347
timestamp 1698431365
transform 1 0 40208 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_6
timestamp 1698431365
transform 1 0 2016 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_42
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_46
timestamp 1698431365
transform 1 0 6496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_50
timestamp 1698431365
transform 1 0 6944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_58
timestamp 1698431365
transform 1 0 7840 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_65
timestamp 1698431365
transform 1 0 8624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_84
timestamp 1698431365
transform 1 0 10752 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_92
timestamp 1698431365
transform 1 0 11648 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_105
timestamp 1698431365
transform 1 0 13104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_109
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_125
timestamp 1698431365
transform 1 0 15344 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_133
timestamp 1698431365
transform 1 0 16240 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_137
timestamp 1698431365
transform 1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_221
timestamp 1698431365
transform 1 0 26096 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_229
timestamp 1698431365
transform 1 0 26992 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_261
timestamp 1698431365
transform 1 0 30576 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_315
timestamp 1698431365
transform 1 0 36624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_319
timestamp 1698431365
transform 1 0 37072 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_335
timestamp 1698431365
transform 1 0 38864 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_343
timestamp 1698431365
transform 1 0 39760 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_347
timestamp 1698431365
transform 1 0 40208 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_43
timestamp 1698431365
transform 1 0 6160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_68
timestamp 1698431365
transform 1 0 8960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_80
timestamp 1698431365
transform 1 0 10304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_84
timestamp 1698431365
transform 1 0 10752 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_100
timestamp 1698431365
transform 1 0 12544 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_119
timestamp 1698431365
transform 1 0 14672 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_125
timestamp 1698431365
transform 1 0 15344 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_133
timestamp 1698431365
transform 1 0 16240 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_152
timestamp 1698431365
transform 1 0 18368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_162
timestamp 1698431365
transform 1 0 19488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_164
timestamp 1698431365
transform 1 0 19712 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_183
timestamp 1698431365
transform 1 0 21840 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_191
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_197
timestamp 1698431365
transform 1 0 23408 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_201
timestamp 1698431365
transform 1 0 23856 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_214
timestamp 1698431365
transform 1 0 25312 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_230
timestamp 1698431365
transform 1 0 27104 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_234
timestamp 1698431365
transform 1 0 27552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_236
timestamp 1698431365
transform 1 0 27776 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_252
timestamp 1698431365
transform 1 0 29568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_268
timestamp 1698431365
transform 1 0 31360 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_272
timestamp 1698431365
transform 1 0 31808 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_275
timestamp 1698431365
transform 1 0 32144 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_279
timestamp 1698431365
transform 1 0 32592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_287
timestamp 1698431365
transform 1 0 33488 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_291
timestamp 1698431365
transform 1 0 33936 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_307
timestamp 1698431365
transform 1 0 35728 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_333
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_341
timestamp 1698431365
transform 1 0 39536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_345
timestamp 1698431365
transform 1 0 39984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_347
timestamp 1698431365
transform 1 0 40208 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_26
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_42
timestamp 1698431365
transform 1 0 6048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_49
timestamp 1698431365
transform 1 0 6832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_65
timestamp 1698431365
transform 1 0 8624 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_84
timestamp 1698431365
transform 1 0 10752 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_86
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_93
timestamp 1698431365
transform 1 0 11760 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_101
timestamp 1698431365
transform 1 0 12656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_105
timestamp 1698431365
transform 1 0 13104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_123
timestamp 1698431365
transform 1 0 15120 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_125
timestamp 1698431365
transform 1 0 15344 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_152
timestamp 1698431365
transform 1 0 18368 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_156
timestamp 1698431365
transform 1 0 18816 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_159
timestamp 1698431365
transform 1 0 19152 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_163
timestamp 1698431365
transform 1 0 19600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_165
timestamp 1698431365
transform 1 0 19824 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_174
timestamp 1698431365
transform 1 0 20832 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_178
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_218
timestamp 1698431365
transform 1 0 25760 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_234
timestamp 1698431365
transform 1 0 27552 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_240
timestamp 1698431365
transform 1 0 28224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_246
timestamp 1698431365
transform 1 0 28896 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_273
timestamp 1698431365
transform 1 0 31920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_294
timestamp 1698431365
transform 1 0 34272 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_326
timestamp 1698431365
transform 1 0 37856 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_342
timestamp 1698431365
transform 1 0 39648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_44
timestamp 1698431365
transform 1 0 6272 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_52
timestamp 1698431365
transform 1 0 7168 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_86
timestamp 1698431365
transform 1 0 10976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_90
timestamp 1698431365
transform 1 0 11424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_96
timestamp 1698431365
transform 1 0 12096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_166
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_201
timestamp 1698431365
transform 1 0 23856 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_209
timestamp 1698431365
transform 1 0 24752 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_213
timestamp 1698431365
transform 1 0 25200 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_233
timestamp 1698431365
transform 1 0 27440 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_251
timestamp 1698431365
transform 1 0 29456 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_253
timestamp 1698431365
transform 1 0 29680 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_321
timestamp 1698431365
transform 1 0 37296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_333
timestamp 1698431365
transform 1 0 38640 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_31
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_35
timestamp 1698431365
transform 1 0 5264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_37
timestamp 1698431365
transform 1 0 5488 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_43
timestamp 1698431365
transform 1 0 6160 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_51
timestamp 1698431365
transform 1 0 7056 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_55
timestamp 1698431365
transform 1 0 7504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_57
timestamp 1698431365
transform 1 0 7728 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_82
timestamp 1698431365
transform 1 0 10528 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_132
timestamp 1698431365
transform 1 0 16128 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_162
timestamp 1698431365
transform 1 0 19488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_166
timestamp 1698431365
transform 1 0 19936 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_170
timestamp 1698431365
transform 1 0 20384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_174
timestamp 1698431365
transform 1 0 20832 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_247
timestamp 1698431365
transform 1 0 29008 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_251
timestamp 1698431365
transform 1 0 29456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_253
timestamp 1698431365
transform 1 0 29680 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_315
timestamp 1698431365
transform 1 0 36624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_319
timestamp 1698431365
transform 1 0 37072 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_335
timestamp 1698431365
transform 1 0 38864 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_343
timestamp 1698431365
transform 1 0 39760 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_18
timestamp 1698431365
transform 1 0 3360 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_26
timestamp 1698431365
transform 1 0 4256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_28
timestamp 1698431365
transform 1 0 4480 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_53
timestamp 1698431365
transform 1 0 7280 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_85
timestamp 1698431365
transform 1 0 10864 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_93
timestamp 1698431365
transform 1 0 11760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_134
timestamp 1698431365
transform 1 0 16352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_140
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_162
timestamp 1698431365
transform 1 0 19488 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_195
timestamp 1698431365
transform 1 0 23184 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_259
timestamp 1698431365
transform 1 0 30352 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_333
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_344
timestamp 1698431365
transform 1 0 39872 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_46
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_50
timestamp 1698431365
transform 1 0 6944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_60
timestamp 1698431365
transform 1 0 8064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_81
timestamp 1698431365
transform 1 0 10416 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_85
timestamp 1698431365
transform 1 0 10864 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_89
timestamp 1698431365
transform 1 0 11312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_96
timestamp 1698431365
transform 1 0 12096 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_108
timestamp 1698431365
transform 1 0 13440 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_119
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_123
timestamp 1698431365
transform 1 0 15120 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_127
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_131
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_144
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_169
timestamp 1698431365
transform 1 0 20272 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_177
timestamp 1698431365
transform 1 0 21168 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_235
timestamp 1698431365
transform 1 0 27664 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_251
timestamp 1698431365
transform 1 0 29456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_253
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_261
timestamp 1698431365
transform 1 0 30576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_272
timestamp 1698431365
transform 1 0 31808 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_288
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_344
timestamp 1698431365
transform 1 0 39872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_62
timestamp 1698431365
transform 1 0 8288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_66
timestamp 1698431365
transform 1 0 8736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_70
timestamp 1698431365
transform 1 0 9184 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_77
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_93
timestamp 1698431365
transform 1 0 11760 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_131
timestamp 1698431365
transform 1 0 16016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_137
timestamp 1698431365
transform 1 0 16688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_139
timestamp 1698431365
transform 1 0 16912 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_142
timestamp 1698431365
transform 1 0 17248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_144
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_153
timestamp 1698431365
transform 1 0 18480 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_155
timestamp 1698431365
transform 1 0 18704 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_162
timestamp 1698431365
transform 1 0 19488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_170
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_181
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_183
timestamp 1698431365
transform 1 0 21840 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_190
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_194
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_199
timestamp 1698431365
transform 1 0 23632 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_203
timestamp 1698431365
transform 1 0 24080 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_210
timestamp 1698431365
transform 1 0 24864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_214
timestamp 1698431365
transform 1 0 25312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_218
timestamp 1698431365
transform 1 0 25760 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_234
timestamp 1698431365
transform 1 0 27552 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_263
timestamp 1698431365
transform 1 0 30800 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_275
timestamp 1698431365
transform 1 0 32144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_283
timestamp 1698431365
transform 1 0 33040 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_300
timestamp 1698431365
transform 1 0 34944 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_308
timestamp 1698431365
transform 1 0 35840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_319
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_344
timestamp 1698431365
transform 1 0 39872 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_22
timestamp 1698431365
transform 1 0 3808 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_32
timestamp 1698431365
transform 1 0 4928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_36
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_47
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_49
timestamp 1698431365
transform 1 0 6832 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698431365
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_104
timestamp 1698431365
transform 1 0 12992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_157
timestamp 1698431365
transform 1 0 18928 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_166
timestamp 1698431365
transform 1 0 19936 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_198
timestamp 1698431365
transform 1 0 23520 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_244
timestamp 1698431365
transform 1 0 28672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_246
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_265
timestamp 1698431365
transform 1 0 31024 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_273
timestamp 1698431365
transform 1 0 31920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_288
timestamp 1698431365
transform 1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_307
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_47
timestamp 1698431365
transform 1 0 6608 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_85
timestamp 1698431365
transform 1 0 10864 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_131
timestamp 1698431365
transform 1 0 16016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_160
timestamp 1698431365
transform 1 0 19264 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_168
timestamp 1698431365
transform 1 0 20160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698431365
transform 1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_193
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_201
timestamp 1698431365
transform 1 0 23856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_205
timestamp 1698431365
transform 1 0 24304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_209
timestamp 1698431365
transform 1 0 24752 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_213
timestamp 1698431365
transform 1 0 25200 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_221
timestamp 1698431365
transform 1 0 26096 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_225
timestamp 1698431365
transform 1 0 26544 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_282
timestamp 1698431365
transform 1 0 32928 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_286
timestamp 1698431365
transform 1 0 33376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_298
timestamp 1698431365
transform 1 0 34720 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_314
timestamp 1698431365
transform 1 0 36512 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_18
timestamp 1698431365
transform 1 0 3360 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_29
timestamp 1698431365
transform 1 0 4592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_33
timestamp 1698431365
transform 1 0 5040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_47
timestamp 1698431365
transform 1 0 6608 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_96
timestamp 1698431365
transform 1 0 12096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_100
timestamp 1698431365
transform 1 0 12544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_108
timestamp 1698431365
transform 1 0 13440 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_116
timestamp 1698431365
transform 1 0 14336 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_132
timestamp 1698431365
transform 1 0 16128 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_149
timestamp 1698431365
transform 1 0 18032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_153
timestamp 1698431365
transform 1 0 18480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_155
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_158
timestamp 1698431365
transform 1 0 19040 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_162
timestamp 1698431365
transform 1 0 19488 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_169
timestamp 1698431365
transform 1 0 20272 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_173
timestamp 1698431365
transform 1 0 20720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_177
timestamp 1698431365
transform 1 0 21168 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_219
timestamp 1698431365
transform 1 0 25872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_221
timestamp 1698431365
transform 1 0 26096 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_308
timestamp 1698431365
transform 1 0 35840 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_317
timestamp 1698431365
transform 1 0 36848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_319
timestamp 1698431365
transform 1 0 37072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_330
timestamp 1698431365
transform 1 0 38304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_344
timestamp 1698431365
transform 1 0 39872 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_12
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_48
timestamp 1698431365
transform 1 0 6720 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_76
timestamp 1698431365
transform 1 0 9856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_80
timestamp 1698431365
transform 1 0 10304 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_89
timestamp 1698431365
transform 1 0 11312 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_93
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_127
timestamp 1698431365
transform 1 0 15568 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_135
timestamp 1698431365
transform 1 0 16464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_139
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_184
timestamp 1698431365
transform 1 0 21952 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_192
timestamp 1698431365
transform 1 0 22848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_196
timestamp 1698431365
transform 1 0 23296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_198
timestamp 1698431365
transform 1 0 23520 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_203
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_249
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_256
timestamp 1698431365
transform 1 0 30016 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_275
timestamp 1698431365
transform 1 0 32144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_277
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_284
timestamp 1698431365
transform 1 0 33152 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_300
timestamp 1698431365
transform 1 0 34944 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_330
timestamp 1698431365
transform 1 0 38304 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_50
timestamp 1698431365
transform 1 0 6944 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_58
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_88
timestamp 1698431365
transform 1 0 11200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_120
timestamp 1698431365
transform 1 0 14784 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_151
timestamp 1698431365
transform 1 0 18256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_155
timestamp 1698431365
transform 1 0 18704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_165
timestamp 1698431365
transform 1 0 19824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_185
timestamp 1698431365
transform 1 0 22064 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_201
timestamp 1698431365
transform 1 0 23856 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_227
timestamp 1698431365
transform 1 0 26768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_229
timestamp 1698431365
transform 1 0 26992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_236
timestamp 1698431365
transform 1 0 27776 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_252
timestamp 1698431365
transform 1 0 29568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_254
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_257
timestamp 1698431365
transform 1 0 30128 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_265
timestamp 1698431365
transform 1 0 31024 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_284
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_306
timestamp 1698431365
transform 1 0 35616 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_329
timestamp 1698431365
transform 1 0 38192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_333
timestamp 1698431365
transform 1 0 38640 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_344
timestamp 1698431365
transform 1 0 39872 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_52
timestamp 1698431365
transform 1 0 7168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_68
timestamp 1698431365
transform 1 0 8960 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_81
timestamp 1698431365
transform 1 0 10416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_85
timestamp 1698431365
transform 1 0 10864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_87
timestamp 1698431365
transform 1 0 11088 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1698431365
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_112
timestamp 1698431365
transform 1 0 13888 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_128
timestamp 1698431365
transform 1 0 15680 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_169
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698431365
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_185
timestamp 1698431365
transform 1 0 22064 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_217
timestamp 1698431365
transform 1 0 25648 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_233
timestamp 1698431365
transform 1 0 27440 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_10
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_12
timestamp 1698431365
transform 1 0 2688 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_24
timestamp 1698431365
transform 1 0 4032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_26
timestamp 1698431365
transform 1 0 4256 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_65
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_114
timestamp 1698431365
transform 1 0 14112 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_146
timestamp 1698431365
transform 1 0 17696 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_163
timestamp 1698431365
transform 1 0 19600 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_171
timestamp 1698431365
transform 1 0 20496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_202
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_223
timestamp 1698431365
transform 1 0 26320 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_227
timestamp 1698431365
transform 1 0 26768 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_230
timestamp 1698431365
transform 1 0 27104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_232
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_241
timestamp 1698431365
transform 1 0 28336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_243
timestamp 1698431365
transform 1 0 28560 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_248
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_255
timestamp 1698431365
transform 1 0 29904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_259
timestamp 1698431365
transform 1 0 30352 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_267
timestamp 1698431365
transform 1 0 31248 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_306
timestamp 1698431365
transform 1 0 35616 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_315
timestamp 1698431365
transform 1 0 36624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_331
timestamp 1698431365
transform 1 0 38416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_333
timestamp 1698431365
transform 1 0 38640 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_39
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_50
timestamp 1698431365
transform 1 0 6944 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_82
timestamp 1698431365
transform 1 0 10528 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_99
timestamp 1698431365
transform 1 0 12432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_142
timestamp 1698431365
transform 1 0 17248 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_146
timestamp 1698431365
transform 1 0 17696 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_153
timestamp 1698431365
transform 1 0 18480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_157
timestamp 1698431365
transform 1 0 18928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_165
timestamp 1698431365
transform 1 0 19824 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_183
timestamp 1698431365
transform 1 0 21840 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_191
timestamp 1698431365
transform 1 0 22736 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_221
timestamp 1698431365
transform 1 0 26096 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_254
timestamp 1698431365
transform 1 0 29792 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_270
timestamp 1698431365
transform 1 0 31584 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_278
timestamp 1698431365
transform 1 0 32480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_299
timestamp 1698431365
transform 1 0 34832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_313
timestamp 1698431365
transform 1 0 36400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_334
timestamp 1698431365
transform 1 0 38752 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_342
timestamp 1698431365
transform 1 0 39648 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_346
timestamp 1698431365
transform 1 0 40096 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_55
timestamp 1698431365
transform 1 0 7504 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_63
timestamp 1698431365
transform 1 0 8400 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_74
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_83
timestamp 1698431365
transform 1 0 10640 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_91
timestamp 1698431365
transform 1 0 11536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_95
timestamp 1698431365
transform 1 0 11984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_151
timestamp 1698431365
transform 1 0 18256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_155
timestamp 1698431365
transform 1 0 18704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_157
timestamp 1698431365
transform 1 0 18928 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_261
timestamp 1698431365
transform 1 0 30576 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_292
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_298
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_306
timestamp 1698431365
transform 1 0 35616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_310
timestamp 1698431365
transform 1 0 36064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_317
timestamp 1698431365
transform 1 0 36848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_319
timestamp 1698431365
transform 1 0 37072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_326
timestamp 1698431365
transform 1 0 37856 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_342
timestamp 1698431365
transform 1 0 39648 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_16
timestamp 1698431365
transform 1 0 3136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_20
timestamp 1698431365
transform 1 0 3584 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_27
timestamp 1698431365
transform 1 0 4368 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_49
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_55
timestamp 1698431365
transform 1 0 7504 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_62
timestamp 1698431365
transform 1 0 8288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_92
timestamp 1698431365
transform 1 0 11648 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_155
timestamp 1698431365
transform 1 0 18704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_159
timestamp 1698431365
transform 1 0 19152 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_161
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_197
timestamp 1698431365
transform 1 0 23408 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_208
timestamp 1698431365
transform 1 0 24640 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_240
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_251
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_287
timestamp 1698431365
transform 1 0 33488 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_303
timestamp 1698431365
transform 1 0 35280 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_37
timestamp 1698431365
transform 1 0 5488 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_41
timestamp 1698431365
transform 1 0 5936 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_60
timestamp 1698431365
transform 1 0 8064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_87
timestamp 1698431365
transform 1 0 11088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_89
timestamp 1698431365
transform 1 0 11312 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_119
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_151
timestamp 1698431365
transform 1 0 18256 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_167
timestamp 1698431365
transform 1 0 20048 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_171
timestamp 1698431365
transform 1 0 20496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_180
timestamp 1698431365
transform 1 0 21504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_182
timestamp 1698431365
transform 1 0 21728 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_189
timestamp 1698431365
transform 1 0 22512 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_205
timestamp 1698431365
transform 1 0 24304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_260
timestamp 1698431365
transform 1 0 30464 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_306
timestamp 1698431365
transform 1 0 35616 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_314
timestamp 1698431365
transform 1 0 36512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_316
timestamp 1698431365
transform 1 0 36736 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_72
timestamp 1698431365
transform 1 0 9408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_74
timestamp 1698431365
transform 1 0 9632 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_88
timestamp 1698431365
transform 1 0 11200 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_92
timestamp 1698431365
transform 1 0 11648 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_100
timestamp 1698431365
transform 1 0 12544 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_136
timestamp 1698431365
transform 1 0 16576 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_152
timestamp 1698431365
transform 1 0 18368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_154
timestamp 1698431365
transform 1 0 18592 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_161
timestamp 1698431365
transform 1 0 19376 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_169
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_173
timestamp 1698431365
transform 1 0 20720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_213
timestamp 1698431365
transform 1 0 25200 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_251
timestamp 1698431365
transform 1 0 29456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_253
timestamp 1698431365
transform 1 0 29680 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_296
timestamp 1698431365
transform 1 0 34496 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_333
timestamp 1698431365
transform 1 0 38640 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_341
timestamp 1698431365
transform 1 0 39536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_345
timestamp 1698431365
transform 1 0 39984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_347
timestamp 1698431365
transform 1 0 40208 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_12
timestamp 1698431365
transform 1 0 2688 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_20
timestamp 1698431365
transform 1 0 3584 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_27
timestamp 1698431365
transform 1 0 4368 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_59
timestamp 1698431365
transform 1 0 7952 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_67
timestamp 1698431365
transform 1 0 8848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698431365
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_162
timestamp 1698431365
transform 1 0 19488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_168
timestamp 1698431365
transform 1 0 20160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_172
timestamp 1698431365
transform 1 0 20608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_177
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_193
timestamp 1698431365
transform 1 0 22960 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_200
timestamp 1698431365
transform 1 0 23744 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_230
timestamp 1698431365
transform 1 0 27104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_232
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_262
timestamp 1698431365
transform 1 0 30688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_266
timestamp 1698431365
transform 1 0 31136 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_292
timestamp 1698431365
transform 1 0 34048 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_296
timestamp 1698431365
transform 1 0 34496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_323
timestamp 1698431365
transform 1 0 37520 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_339
timestamp 1698431365
transform 1 0 39312 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_41
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_48
timestamp 1698431365
transform 1 0 6720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_52
timestamp 1698431365
transform 1 0 7168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_68
timestamp 1698431365
transform 1 0 8960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_76
timestamp 1698431365
transform 1 0 9856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_80
timestamp 1698431365
transform 1 0 10304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_84
timestamp 1698431365
transform 1 0 10752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_88
timestamp 1698431365
transform 1 0 11200 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_92
timestamp 1698431365
transform 1 0 11648 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_123
timestamp 1698431365
transform 1 0 15120 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_127
timestamp 1698431365
transform 1 0 15568 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_156
timestamp 1698431365
transform 1 0 18816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_166
timestamp 1698431365
transform 1 0 19936 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_206
timestamp 1698431365
transform 1 0 24416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_210
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_214
timestamp 1698431365
transform 1 0 25312 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_240
timestamp 1698431365
transform 1 0 28224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_258
timestamp 1698431365
transform 1 0 30240 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_266
timestamp 1698431365
transform 1 0 31136 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_287
timestamp 1698431365
transform 1 0 33488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_289
timestamp 1698431365
transform 1 0 33712 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_338
timestamp 1698431365
transform 1 0 39200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_57
timestamp 1698431365
transform 1 0 7728 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_65
timestamp 1698431365
transform 1 0 8624 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698431365
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_132
timestamp 1698431365
transform 1 0 16128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_159
timestamp 1698431365
transform 1 0 19152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_163
timestamp 1698431365
transform 1 0 19600 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_179
timestamp 1698431365
transform 1 0 21392 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_187
timestamp 1698431365
transform 1 0 22288 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_194
timestamp 1698431365
transform 1 0 23072 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_216
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_228
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_242
timestamp 1698431365
transform 1 0 28448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_258
timestamp 1698431365
transform 1 0 30240 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_266
timestamp 1698431365
transform 1 0 31136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_270
timestamp 1698431365
transform 1 0 31584 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_278
timestamp 1698431365
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_289
timestamp 1698431365
transform 1 0 33712 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_297
timestamp 1698431365
transform 1 0 34608 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_301
timestamp 1698431365
transform 1 0 35056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_315
timestamp 1698431365
transform 1 0 36624 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_347
timestamp 1698431365
transform 1 0 40208 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_84
timestamp 1698431365
transform 1 0 10752 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_130
timestamp 1698431365
transform 1 0 15904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_134
timestamp 1698431365
transform 1 0 16352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_168
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_185
timestamp 1698431365
transform 1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_187
timestamp 1698431365
transform 1 0 22288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_190
timestamp 1698431365
transform 1 0 22624 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_198
timestamp 1698431365
transform 1 0 23520 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_207
timestamp 1698431365
transform 1 0 24528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_240
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_259
timestamp 1698431365
transform 1 0 30352 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_273
timestamp 1698431365
transform 1 0 31920 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_289
timestamp 1698431365
transform 1 0 33712 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_297
timestamp 1698431365
transform 1 0 34608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_301
timestamp 1698431365
transform 1 0 35056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_308
timestamp 1698431365
transform 1 0 35840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698431365
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_327
timestamp 1698431365
transform 1 0 37968 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_334
timestamp 1698431365
transform 1 0 38752 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_342
timestamp 1698431365
transform 1 0 39648 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_346
timestamp 1698431365
transform 1 0 40096 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_34
timestamp 1698431365
transform 1 0 5152 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_50
timestamp 1698431365
transform 1 0 6944 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_82
timestamp 1698431365
transform 1 0 10528 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_112
timestamp 1698431365
transform 1 0 13888 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_116
timestamp 1698431365
transform 1 0 14336 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_119
timestamp 1698431365
transform 1 0 14672 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_147
timestamp 1698431365
transform 1 0 17808 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_188
timestamp 1698431365
transform 1 0 22400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_231
timestamp 1698431365
transform 1 0 27216 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_247
timestamp 1698431365
transform 1 0 29008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_249
timestamp 1698431365
transform 1 0 29232 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_255
timestamp 1698431365
transform 1 0 29904 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_259
timestamp 1698431365
transform 1 0 30352 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_266
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_270
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_275
timestamp 1698431365
transform 1 0 32144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_292
timestamp 1698431365
transform 1 0 34048 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_300
timestamp 1698431365
transform 1 0 34944 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_304
timestamp 1698431365
transform 1 0 35392 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_312
timestamp 1698431365
transform 1 0 36288 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_316
timestamp 1698431365
transform 1 0 36736 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_66
timestamp 1698431365
transform 1 0 8736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_83
timestamp 1698431365
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_87
timestamp 1698431365
transform 1 0 11088 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_95
timestamp 1698431365
transform 1 0 11984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_99
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_139
timestamp 1698431365
transform 1 0 16912 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_143
timestamp 1698431365
transform 1 0 17360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_161
timestamp 1698431365
transform 1 0 19376 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_169
timestamp 1698431365
transform 1 0 20272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_179
timestamp 1698431365
transform 1 0 21392 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_198
timestamp 1698431365
transform 1 0 23520 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_214
timestamp 1698431365
transform 1 0 25312 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_226
timestamp 1698431365
transform 1 0 26656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_253
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_284
timestamp 1698431365
transform 1 0 33152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_286
timestamp 1698431365
transform 1 0 33376 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_299
timestamp 1698431365
transform 1 0 34832 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_307
timestamp 1698431365
transform 1 0 35728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_333
timestamp 1698431365
transform 1 0 38640 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_341
timestamp 1698431365
transform 1 0 39536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_345
timestamp 1698431365
transform 1 0 39984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_347
timestamp 1698431365
transform 1 0 40208 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_80
timestamp 1698431365
transform 1 0 10304 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_94
timestamp 1698431365
transform 1 0 11872 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_124
timestamp 1698431365
transform 1 0 15232 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_146
timestamp 1698431365
transform 1 0 17696 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_154
timestamp 1698431365
transform 1 0 18592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_161
timestamp 1698431365
transform 1 0 19376 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_193
timestamp 1698431365
transform 1 0 22960 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_197
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_207
timestamp 1698431365
transform 1 0 24528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_214
timestamp 1698431365
transform 1 0 25312 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_228
timestamp 1698431365
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_298
timestamp 1698431365
transform 1 0 34720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_317
timestamp 1698431365
transform 1 0 36848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_53
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_63
timestamp 1698431365
transform 1 0 8400 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_67
timestamp 1698431365
transform 1 0 8848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_72
timestamp 1698431365
transform 1 0 9408 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_88
timestamp 1698431365
transform 1 0 11200 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_96
timestamp 1698431365
transform 1 0 12096 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_138
timestamp 1698431365
transform 1 0 16800 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_146
timestamp 1698431365
transform 1 0 17696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_148
timestamp 1698431365
transform 1 0 17920 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_161
timestamp 1698431365
transform 1 0 19376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_163
timestamp 1698431365
transform 1 0 19600 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_188
timestamp 1698431365
transform 1 0 22400 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_192
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_216
timestamp 1698431365
transform 1 0 25536 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_218
timestamp 1698431365
transform 1 0 25760 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_221
timestamp 1698431365
transform 1 0 26096 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_223
timestamp 1698431365
transform 1 0 26320 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_300
timestamp 1698431365
transform 1 0 34944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_331
timestamp 1698431365
transform 1 0 38416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_335
timestamp 1698431365
transform 1 0 38864 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_343
timestamp 1698431365
transform 1 0 39760 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_347
timestamp 1698431365
transform 1 0 40208 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_34
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_50
timestamp 1698431365
transform 1 0 6944 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_54
timestamp 1698431365
transform 1 0 7392 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_84
timestamp 1698431365
transform 1 0 10752 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_138
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_148
timestamp 1698431365
transform 1 0 17920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_152
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_181
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_197
timestamp 1698431365
transform 1 0 23408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_201
timestamp 1698431365
transform 1 0 23856 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_214
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_223
timestamp 1698431365
transform 1 0 26320 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_227
timestamp 1698431365
transform 1 0 26768 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_230
timestamp 1698431365
transform 1 0 27104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_234
timestamp 1698431365
transform 1 0 27552 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_242
timestamp 1698431365
transform 1 0 28448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_244
timestamp 1698431365
transform 1 0 28672 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_327
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_343
timestamp 1698431365
transform 1 0 39760 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_347
timestamp 1698431365
transform 1 0 40208 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_78
timestamp 1698431365
transform 1 0 10080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_80
timestamp 1698431365
transform 1 0 10304 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_94
timestamp 1698431365
transform 1 0 11872 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_113
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_136
timestamp 1698431365
transform 1 0 16576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_140
timestamp 1698431365
transform 1 0 17024 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_148
timestamp 1698431365
transform 1 0 17920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_150
timestamp 1698431365
transform 1 0 18144 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_169
timestamp 1698431365
transform 1 0 20272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_173
timestamp 1698431365
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_181
timestamp 1698431365
transform 1 0 21616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_183
timestamp 1698431365
transform 1 0 21840 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_190
timestamp 1698431365
transform 1 0 22624 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_206
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_239
timestamp 1698431365
transform 1 0 28112 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_278
timestamp 1698431365
transform 1 0 32480 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_294
timestamp 1698431365
transform 1 0 34272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_298
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_337
timestamp 1698431365
transform 1 0 39088 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_345
timestamp 1698431365
transform 1 0 39984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_347
timestamp 1698431365
transform 1 0 40208 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_34
timestamp 1698431365
transform 1 0 5152 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_50
timestamp 1698431365
transform 1 0 6944 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_54
timestamp 1698431365
transform 1 0 7392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_62
timestamp 1698431365
transform 1 0 8288 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_100
timestamp 1698431365
transform 1 0 12544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_104
timestamp 1698431365
transform 1 0 12992 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_111
timestamp 1698431365
transform 1 0 13776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_113
timestamp 1698431365
transform 1 0 14000 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_116
timestamp 1698431365
transform 1 0 14336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_164
timestamp 1698431365
transform 1 0 19712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_174
timestamp 1698431365
transform 1 0 20832 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_190
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_194
timestamp 1698431365
transform 1 0 23072 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_196
timestamp 1698431365
transform 1 0 23296 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_207
timestamp 1698431365
transform 1 0 24528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_216
timestamp 1698431365
transform 1 0 25536 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_223
timestamp 1698431365
transform 1 0 26320 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_239
timestamp 1698431365
transform 1 0 28112 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_255
timestamp 1698431365
transform 1 0 29904 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_261
timestamp 1698431365
transform 1 0 30576 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_270
timestamp 1698431365
transform 1 0 31584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_274
timestamp 1698431365
transform 1 0 32032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_278
timestamp 1698431365
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_294
timestamp 1698431365
transform 1 0 34272 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_326
timestamp 1698431365
transform 1 0 37856 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_342
timestamp 1698431365
transform 1 0 39648 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_69
timestamp 1698431365
transform 1 0 9072 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_97
timestamp 1698431365
transform 1 0 12208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_115
timestamp 1698431365
transform 1 0 14224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_117
timestamp 1698431365
transform 1 0 14448 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_127
timestamp 1698431365
transform 1 0 15568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_131
timestamp 1698431365
transform 1 0 16016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_133
timestamp 1698431365
transform 1 0 16240 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_136
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_140
timestamp 1698431365
transform 1 0 17024 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_148
timestamp 1698431365
transform 1 0 17920 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_152
timestamp 1698431365
transform 1 0 18368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_154
timestamp 1698431365
transform 1 0 18592 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_165
timestamp 1698431365
transform 1 0 19824 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_189
timestamp 1698431365
transform 1 0 22512 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_191
timestamp 1698431365
transform 1 0 22736 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_229
timestamp 1698431365
transform 1 0 26992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_233
timestamp 1698431365
transform 1 0 27440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_298
timestamp 1698431365
transform 1 0 34720 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698431365
transform 1 0 38640 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_341
timestamp 1698431365
transform 1 0 39536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_345
timestamp 1698431365
transform 1 0 39984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_347
timestamp 1698431365
transform 1 0 40208 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_50
timestamp 1698431365
transform 1 0 6944 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_58
timestamp 1698431365
transform 1 0 7840 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_65
timestamp 1698431365
transform 1 0 8624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_97
timestamp 1698431365
transform 1 0 12208 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_105
timestamp 1698431365
transform 1 0 13104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_115
timestamp 1698431365
transform 1 0 14224 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_123
timestamp 1698431365
transform 1 0 15120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_125
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_131
timestamp 1698431365
transform 1 0 16016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_147
timestamp 1698431365
transform 1 0 17808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_151
timestamp 1698431365
transform 1 0 18256 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_167
timestamp 1698431365
transform 1 0 20048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_169
timestamp 1698431365
transform 1 0 20272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_176
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_192
timestamp 1698431365
transform 1 0 22848 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_201
timestamp 1698431365
transform 1 0 23856 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_205
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_207
timestamp 1698431365
transform 1 0 24528 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_318
timestamp 1698431365
transform 1 0 36960 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_334
timestamp 1698431365
transform 1 0 38752 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_342
timestamp 1698431365
transform 1 0 39648 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_6
timestamp 1698431365
transform 1 0 2016 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_22
timestamp 1698431365
transform 1 0 3808 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_30
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_82
timestamp 1698431365
transform 1 0 10528 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_90
timestamp 1698431365
transform 1 0 11424 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_103
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_116
timestamp 1698431365
transform 1 0 14336 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_125
timestamp 1698431365
transform 1 0 15344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_127
timestamp 1698431365
transform 1 0 15568 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_186
timestamp 1698431365
transform 1 0 22176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_188
timestamp 1698431365
transform 1 0 22400 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_191
timestamp 1698431365
transform 1 0 22736 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_207
timestamp 1698431365
transform 1 0 24528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_221
timestamp 1698431365
transform 1 0 26096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_231
timestamp 1698431365
transform 1 0 27216 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_239
timestamp 1698431365
transform 1 0 28112 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_253
timestamp 1698431365
transform 1 0 29680 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_261
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_265
timestamp 1698431365
transform 1 0 31024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_269
timestamp 1698431365
transform 1 0 31472 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_301
timestamp 1698431365
transform 1 0 35056 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_309
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_333
timestamp 1698431365
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_341
timestamp 1698431365
transform 1 0 39536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_345
timestamp 1698431365
transform 1 0 39984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_347
timestamp 1698431365
transform 1 0 40208 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_6
timestamp 1698431365
transform 1 0 2016 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_78
timestamp 1698431365
transform 1 0 10080 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_94
timestamp 1698431365
transform 1 0 11872 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_102
timestamp 1698431365
transform 1 0 12768 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_115
timestamp 1698431365
transform 1 0 14224 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_149
timestamp 1698431365
transform 1 0 18032 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_157
timestamp 1698431365
transform 1 0 18928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_161
timestamp 1698431365
transform 1 0 19376 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_197
timestamp 1698431365
transform 1 0 23408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698431365
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_222
timestamp 1698431365
transform 1 0 26208 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_236
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_240
timestamp 1698431365
transform 1 0 28224 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_256
timestamp 1698431365
transform 1 0 30016 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_330
timestamp 1698431365
transform 1 0 38304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_338
timestamp 1698431365
transform 1 0 39200 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_342
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_85
timestamp 1698431365
transform 1 0 10864 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_93
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_103
timestamp 1698431365
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_130
timestamp 1698431365
transform 1 0 15904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_161
timestamp 1698431365
transform 1 0 19376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_165
timestamp 1698431365
transform 1 0 19824 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_183
timestamp 1698431365
transform 1 0 21840 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_199
timestamp 1698431365
transform 1 0 23632 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_228
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_234
timestamp 1698431365
transform 1 0 27552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_280
timestamp 1698431365
transform 1 0 32704 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_312
timestamp 1698431365
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698431365
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_341
timestamp 1698431365
transform 1 0 39536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_343
timestamp 1698431365
transform 1 0 39760 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_84
timestamp 1698431365
transform 1 0 10752 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_86
timestamp 1698431365
transform 1 0 10976 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_116
timestamp 1698431365
transform 1 0 14336 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_132
timestamp 1698431365
transform 1 0 16128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_218
timestamp 1698431365
transform 1 0 25760 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_234
timestamp 1698431365
transform 1 0 27552 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_247
timestamp 1698431365
transform 1 0 29008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_249
timestamp 1698431365
transform 1 0 29232 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_288
timestamp 1698431365
transform 1 0 33600 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_320
timestamp 1698431365
transform 1 0 37184 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_336
timestamp 1698431365
transform 1 0 38976 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_193
timestamp 1698431365
transform 1 0 22960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_195
timestamp 1698431365
transform 1 0 23184 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_225
timestamp 1698431365
transform 1 0 26544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_229
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_236
timestamp 1698431365
transform 1 0 27776 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_253
timestamp 1698431365
transform 1 0 29680 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_283
timestamp 1698431365
transform 1 0 33040 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_333
timestamp 1698431365
transform 1 0 38640 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_341
timestamp 1698431365
transform 1 0 39536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_343
timestamp 1698431365
transform 1 0 39760 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_246
timestamp 1698431365
transform 1 0 28896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_250
timestamp 1698431365
transform 1 0 29344 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_314
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_330
timestamp 1698431365
transform 1 0 38304 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_338
timestamp 1698431365
transform 1 0 39200 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_342
timestamp 1698431365
transform 1 0 39648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_6
timestamp 1698431365
transform 1 0 2016 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_22
timestamp 1698431365
transform 1 0 3808 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_30
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_251
timestamp 1698431365
transform 1 0 29456 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_255
timestamp 1698431365
transform 1 0 29904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_257
timestamp 1698431365
transform 1 0 30128 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_260
timestamp 1698431365
transform 1 0 30464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_264
timestamp 1698431365
transform 1 0 30912 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_296
timestamp 1698431365
transform 1 0 34496 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698431365
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_333
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_337
timestamp 1698431365
transform 1 0 39088 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_339
timestamp 1698431365
transform 1 0 39312 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_36
timestamp 1698431365
transform 1 0 5376 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_52
timestamp 1698431365
transform 1 0 7168 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_60
timestamp 1698431365
transform 1 0 8064 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_65
timestamp 1698431365
transform 1 0 8624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_67
timestamp 1698431365
transform 1 0 8848 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_70
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_240
timestamp 1698431365
transform 1 0 28224 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_312
timestamp 1698431365
transform 1 0 36288 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_328
timestamp 1698431365
transform 1 0 38080 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_342
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 40320 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform -1 0 40320 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 40320 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output8 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output9 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38752 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output10
timestamp 1698431365
transform 1 0 38752 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output11
timestamp 1698431365
transform 1 0 38752 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output12
timestamp 1698431365
transform 1 0 38752 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output13
timestamp 1698431365
transform 1 0 38752 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output14
timestamp 1698431365
transform 1 0 38752 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output15
timestamp 1698431365
transform 1 0 37184 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output16
timestamp 1698431365
transform 1 0 38752 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output17
timestamp 1698431365
transform 1 0 38752 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output18 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1698431365
transform 1 0 38752 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output20
timestamp 1698431365
transform -1 0 3136 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output21
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_50 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_51
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_52
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 40544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_53
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_54
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 40544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_55
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_56
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 40544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_57
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_58
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 40544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_59
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_60
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 40544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_61
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_62
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 40544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 40544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 40544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 40544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 40544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 40544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 40544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 40544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 40544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 40544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 40544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 40544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 40544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 40544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 40544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 40544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 40544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 40544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_28 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39872 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_29
timestamp 1698431365
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_30
timestamp 1698431365
transform 1 0 39424 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_31
timestamp 1698431365
transform -1 0 36288 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_32
timestamp 1698431365
transform -1 0 11312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_33
timestamp 1698431365
transform -1 0 2016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_34
timestamp 1698431365
transform 1 0 39872 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_35
timestamp 1698431365
transform 1 0 39872 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_36
timestamp 1698431365
transform -1 0 10640 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_37
timestamp 1698431365
transform 1 0 38976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_38
timestamp 1698431365
transform -1 0 2016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_39
timestamp 1698431365
transform -1 0 2016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_40
timestamp 1698431365
transform 1 0 39872 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_41
timestamp 1698431365
transform 1 0 39872 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_42
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_43
timestamp 1698431365
transform 1 0 39872 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_44
timestamp 1698431365
transform 1 0 39872 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_45
timestamp 1698431365
transform 1 0 39424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_46
timestamp 1698431365
transform -1 0 8624 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_47
timestamp 1698431365
transform -1 0 2016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_48
timestamp 1698431365
transform -1 0 2016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_49
timestamp 1698431365
transform 1 0 39872 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_50
timestamp 1698431365
transform 1 0 39872 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_51
timestamp 1698431365
transform -1 0 2016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_52
timestamp 1698431365
transform 1 0 39872 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_53
timestamp 1698431365
transform 1 0 38976 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_54
timestamp 1698431365
transform -1 0 2016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_55
timestamp 1698431365
transform 1 0 39872 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_56
timestamp 1698431365
transform 1 0 38528 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_57
timestamp 1698431365
transform -1 0 2016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_58
timestamp 1698431365
transform 1 0 39424 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  solo_squash_caravel_gf180_59
timestamp 1698431365
transform 1 0 39872 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_100 asic_tools/pdk/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_110
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_114
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_115
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_119
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_120
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_121
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_123
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_124
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_125
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_126
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_128
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_129
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_130
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_131
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_132
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_133
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_134
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_135
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_136
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_137
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_138
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_139
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_140
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_141
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_142
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_143
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_144
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_145
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_146
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_147
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_148
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_149
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_150
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_151
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_152
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_153
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_154
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_155
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_156
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_157
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_158
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_159
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_160
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_161
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_162
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_163
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_164
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_165
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_166
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_167
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_168
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_169
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_170
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_171
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_172
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_173
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_174
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_175
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_176
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_177
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_178
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_179
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_180
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_181
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_182
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_183
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_184
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_185
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_186
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_187
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_188
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_189
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_190
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_191
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_192
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_193
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_194
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_195
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_196
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_197
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_198
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_199
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_200
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_201
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_202
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_203
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_204
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_205
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_206
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_207
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_208
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_209
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_210
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_211
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_212
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_213
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_214
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_215
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_216
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_217
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_218
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_219
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_220
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_221
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_222
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_223
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_224
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_225
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_226
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_227
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_228
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_229
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_230
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_231
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_232
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_233
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_234
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_235
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_236
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_237
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_238
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_239
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_240
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_241
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_242
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_243
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_244
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_245
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_246
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_247
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_248
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_249
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_250
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_251
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_252
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_253
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_254
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_255
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_256
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_257
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_258
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_259
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_260
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_261
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_262
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_263
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_264
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_265
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_266
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_267
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_268
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_269
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_270
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_271
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_272
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_273
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_274
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_275
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_276
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_277
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_278
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_279
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_280
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_281
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_282
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_283
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_284
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_285
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_286
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_287
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_288
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_289
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_290
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_291
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_292
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_293
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_294
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_295
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_296
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_297
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_298
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_299
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_300
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_301
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_302
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_303
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_304
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_305
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_306
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_307
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_308
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_309
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_310
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_311
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_312
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_313
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_314
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_315
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_316
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_317
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_318
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_319
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_320
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_321
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_322
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_323
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_324
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_325
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_326
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_327
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_328
timestamp 1698431365
transform 1 0 12768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_329
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_330
timestamp 1698431365
transform 1 0 20384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_331
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_332
timestamp 1698431365
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_333
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_334
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_335
timestamp 1698431365
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
<< labels >>
flabel metal3 s 41101 14784 41901 14896 0 FreeSans 448 0 0 0 blue
port 0 nsew signal tristate
flabel metal3 s 41101 12768 41901 12880 0 FreeSans 448 0 0 0 debug_design_reset
port 1 nsew signal tristate
flabel metal3 s 41101 7392 41901 7504 0 FreeSans 448 0 0 0 debug_gpio_ready
port 2 nsew signal tristate
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 down_key_n
port 3 nsew signal input
flabel metal3 s 41101 26208 41901 26320 0 FreeSans 448 0 0 0 ext_reset_n
port 4 nsew signal input
flabel metal3 s 41101 5376 41901 5488 0 FreeSans 448 0 0 0 gpio_ready
port 5 nsew signal input
flabel metal3 s 41101 20832 41901 20944 0 FreeSans 448 0 0 0 green
port 6 nsew signal tristate
flabel metal3 s 41101 20160 41901 20272 0 FreeSans 448 0 0 0 hsync
port 7 nsew signal tristate
flabel metal3 s 41101 36960 41901 37072 0 FreeSans 448 0 0 0 io_oeb[0]
port 8 nsew signal tristate
flabel metal3 s 0 6048 800 6160 0 FreeSans 448 0 0 0 io_oeb[10]
port 9 nsew signal tristate
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 io_oeb[11]
port 10 nsew signal tristate
flabel metal3 s 41101 40320 41901 40432 0 FreeSans 448 0 0 0 io_oeb[12]
port 11 nsew signal tristate
flabel metal3 s 41101 15456 41901 15568 0 FreeSans 448 0 0 0 io_oeb[13]
port 12 nsew signal tristate
flabel metal3 s 41101 17472 41901 17584 0 FreeSans 448 0 0 0 io_oeb[14]
port 13 nsew signal tristate
flabel metal3 s 41101 18144 41901 18256 0 FreeSans 448 0 0 0 io_oeb[15]
port 14 nsew signal tristate
flabel metal3 s 41101 16800 41901 16912 0 FreeSans 448 0 0 0 io_oeb[16]
port 15 nsew signal tristate
flabel metal3 s 41101 18816 41901 18928 0 FreeSans 448 0 0 0 io_oeb[17]
port 16 nsew signal tristate
flabel metal3 s 41101 16128 41901 16240 0 FreeSans 448 0 0 0 io_oeb[18]
port 17 nsew signal tristate
flabel metal3 s 41101 12096 41901 12208 0 FreeSans 448 0 0 0 io_oeb[19]
port 18 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 19 nsew signal tristate
flabel metal3 s 41101 42336 41901 42448 0 FreeSans 448 0 0 0 io_oeb[20]
port 20 nsew signal tristate
flabel metal3 s 41101 8064 41901 8176 0 FreeSans 448 0 0 0 io_oeb[21]
port 21 nsew signal tristate
flabel metal3 s 41101 39648 41901 39760 0 FreeSans 448 0 0 0 io_oeb[22]
port 22 nsew signal tristate
flabel metal3 s 41101 2688 41901 2800 0 FreeSans 448 0 0 0 io_oeb[23]
port 23 nsew signal tristate
flabel metal2 s 8064 44685 8176 45485 0 FreeSans 448 90 0 0 io_oeb[24]
port 24 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 io_oeb[25]
port 25 nsew signal tristate
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 io_oeb[26]
port 26 nsew signal tristate
flabel metal3 s 41101 38304 41901 38416 0 FreeSans 448 0 0 0 io_oeb[27]
port 27 nsew signal tristate
flabel metal3 s 41101 6048 41901 6160 0 FreeSans 448 0 0 0 io_oeb[28]
port 28 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 io_oeb[29]
port 29 nsew signal tristate
flabel metal3 s 41101 40992 41901 41104 0 FreeSans 448 0 0 0 io_oeb[2]
port 30 nsew signal tristate
flabel metal3 s 41101 37632 41901 37744 0 FreeSans 448 0 0 0 io_oeb[30]
port 31 nsew signal tristate
flabel metal3 s 41101 41664 41901 41776 0 FreeSans 448 0 0 0 io_oeb[31]
port 32 nsew signal tristate
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 io_oeb[32]
port 33 nsew signal tristate
flabel metal3 s 41101 38976 41901 39088 0 FreeSans 448 0 0 0 io_oeb[33]
port 34 nsew signal tristate
flabel metal3 s 41101 43008 41901 43120 0 FreeSans 448 0 0 0 io_oeb[34]
port 35 nsew signal tristate
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 io_oeb[35]
port 36 nsew signal tristate
flabel metal3 s 41101 6720 41901 6832 0 FreeSans 448 0 0 0 io_oeb[36]
port 37 nsew signal tristate
flabel metal3 s 41101 3360 41901 3472 0 FreeSans 448 0 0 0 io_oeb[37]
port 38 nsew signal tristate
flabel metal2 s 35616 44685 35728 45485 0 FreeSans 448 90 0 0 io_oeb[3]
port 39 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 io_oeb[4]
port 40 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 io_oeb[5]
port 41 nsew signal tristate
flabel metal3 s 41101 4704 41901 4816 0 FreeSans 448 0 0 0 io_oeb[6]
port 42 nsew signal tristate
flabel metal3 s 41101 4032 41901 4144 0 FreeSans 448 0 0 0 io_oeb[7]
port 43 nsew signal tristate
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 io_oeb[8]
port 44 nsew signal tristate
flabel metal3 s 41101 2016 41901 2128 0 FreeSans 448 0 0 0 io_oeb[9]
port 45 nsew signal tristate
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 new_game_n
port 46 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 pause_n
port 47 nsew signal input
flabel metal3 s 41101 19488 41901 19600 0 FreeSans 448 0 0 0 red
port 48 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 speaker
port 49 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 up_key_n
port 50 nsew signal input
flabel metal4 s 4448 3076 4768 42396 0 FreeSans 1280 90 0 0 vdd
port 51 nsew power bidirectional
flabel metal4 s 35168 3076 35488 42396 0 FreeSans 1280 90 0 0 vdd
port 51 nsew power bidirectional
flabel metal4 s 19808 3076 20128 42396 0 FreeSans 1280 90 0 0 vss
port 52 nsew ground bidirectional
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 vsync
port 53 nsew signal tristate
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 wb_clk_i
port 54 nsew signal input
flabel metal3 s 41101 26880 41901 26992 0 FreeSans 448 0 0 0 wb_rst_i
port 55 nsew signal input
rlabel metal1 20944 41552 20944 41552 0 vdd
rlabel metal1 20944 42336 20944 42336 0 vss
rlabel metal2 14056 7560 14056 7560 0 _0000_
rlabel metal2 19544 7112 19544 7112 0 _0001_
rlabel metal2 20216 4536 20216 4536 0 _0002_
rlabel metal2 24024 4592 24024 4592 0 _0003_
rlabel metal2 26264 6440 26264 6440 0 _0004_
rlabel metal2 11704 9352 11704 9352 0 _0005_
rlabel metal3 2940 13832 2940 13832 0 _0006_
rlabel metal3 6608 10584 6608 10584 0 _0007_
rlabel metal2 2744 11032 2744 11032 0 _0008_
rlabel metal2 8848 8344 8848 8344 0 _0009_
rlabel metal2 2520 16408 2520 16408 0 _0010_
rlabel metal2 10752 24024 10752 24024 0 _0011_
rlabel metal2 3864 24360 3864 24360 0 _0012_
rlabel metal2 3864 25816 3864 25816 0 _0013_
rlabel metal2 7112 29008 7112 29008 0 _0014_
rlabel metal2 5432 28336 5432 28336 0 _0015_
rlabel metal2 7784 33656 7784 33656 0 _0016_
rlabel metal2 8232 36792 8232 36792 0 _0017_
rlabel metal2 12208 38696 12208 38696 0 _0018_
rlabel metal2 17752 36904 17752 36904 0 _0019_
rlabel metal2 12936 32256 12936 32256 0 _0020_
rlabel metal2 21784 37744 21784 37744 0 _0021_
rlabel metal2 23912 34552 23912 34552 0 _0022_
rlabel metal2 25368 39256 25368 39256 0 _0023_
rlabel metal2 27272 40040 27272 40040 0 _0024_
rlabel metal2 31976 39984 31976 39984 0 _0025_
rlabel metal3 31864 34328 31864 34328 0 _0026_
rlabel metal2 25760 32760 25760 32760 0 _0027_
rlabel metal2 38024 31304 38024 31304 0 _0028_
rlabel metal2 38024 29904 38024 29904 0 _0029_
rlabel metal2 25928 29344 25928 29344 0 _0030_
rlabel metal2 25144 22568 25144 22568 0 _0031_
rlabel metal2 28392 26600 28392 26600 0 _0032_
rlabel metal2 13944 28952 13944 28952 0 _0033_
rlabel metal2 27384 22736 27384 22736 0 _0034_
rlabel metal3 22120 26936 22120 26936 0 _0035_
rlabel metal2 34104 10192 34104 10192 0 _0036_
rlabel metal2 35224 9520 35224 9520 0 _0037_
rlabel metal2 31752 9744 31752 9744 0 _0038_
rlabel metal2 34104 12544 34104 12544 0 _0039_
rlabel metal3 35168 13832 35168 13832 0 _0040_
rlabel metal3 37352 16968 37352 16968 0 _0041_
rlabel metal2 37800 18144 37800 18144 0 _0042_
rlabel metal2 37576 22400 37576 22400 0 _0043_
rlabel metal2 38024 19992 38024 19992 0 _0044_
rlabel metal2 37576 23968 37576 23968 0 _0045_
rlabel metal2 25704 18704 25704 18704 0 _0046_
rlabel metal2 16072 10528 16072 10528 0 _0047_
rlabel metal2 20664 9240 20664 9240 0 _0048_
rlabel metal2 17080 9296 17080 9296 0 _0049_
rlabel metal2 22512 15400 22512 15400 0 _0050_
rlabel metal2 15512 17192 15512 17192 0 _0051_
rlabel metal3 15008 24584 15008 24584 0 _0052_
rlabel metal2 18088 23520 18088 23520 0 _0053_
rlabel metal3 14672 23128 14672 23128 0 _0054_
rlabel metal2 21896 21224 21896 21224 0 _0055_
rlabel metal2 22008 18424 22008 18424 0 _0056_
rlabel metal2 24416 25704 24416 25704 0 _0057_
rlabel metal2 23912 25816 23912 25816 0 _0058_
rlabel metal3 23296 25368 23296 25368 0 _0059_
rlabel metal2 22344 23800 22344 23800 0 _0060_
rlabel metal2 21672 20664 21672 20664 0 _0061_
rlabel metal2 17864 21448 17864 21448 0 _0062_
rlabel metal3 18704 21560 18704 21560 0 _0063_
rlabel metal2 15568 26880 15568 26880 0 _0064_
rlabel metal2 18088 21056 18088 21056 0 _0065_
rlabel metal3 18200 20160 18200 20160 0 _0066_
rlabel metal2 31920 21336 31920 21336 0 _0067_
rlabel metal2 35896 21952 35896 21952 0 _0068_
rlabel metal3 37520 23352 37520 23352 0 _0069_
rlabel metal2 37016 19992 37016 19992 0 _0070_
rlabel metal2 35560 22288 35560 22288 0 _0071_
rlabel metal2 27048 19824 27048 19824 0 _0072_
rlabel metal2 26432 18536 26432 18536 0 _0073_
rlabel metal2 33992 17696 33992 17696 0 _0074_
rlabel metal2 29848 22736 29848 22736 0 _0075_
rlabel metal2 17584 16968 17584 16968 0 _0076_
rlabel metal2 19432 21952 19432 21952 0 _0077_
rlabel metal2 18424 20272 18424 20272 0 _0078_
rlabel metal2 18816 21336 18816 21336 0 _0079_
rlabel metal2 28168 22064 28168 22064 0 _0080_
rlabel metal2 20160 15512 20160 15512 0 _0081_
rlabel metal3 23296 14504 23296 14504 0 _0082_
rlabel metal2 17640 16240 17640 16240 0 _0083_
rlabel metal2 27160 9184 27160 9184 0 _0084_
rlabel metal3 17080 14392 17080 14392 0 _0085_
rlabel metal2 15176 11760 15176 11760 0 _0086_
rlabel metal2 16856 13776 16856 13776 0 _0087_
rlabel metal2 17808 14616 17808 14616 0 _0088_
rlabel metal2 19712 17640 19712 17640 0 _0089_
rlabel metal2 18368 18424 18368 18424 0 _0090_
rlabel metal2 19208 14504 19208 14504 0 _0091_
rlabel metal2 17976 15792 17976 15792 0 _0092_
rlabel metal2 16072 15120 16072 15120 0 _0093_
rlabel metal3 17136 14280 17136 14280 0 _0094_
rlabel metal2 20104 11704 20104 11704 0 _0095_
rlabel metal3 18312 15400 18312 15400 0 _0096_
rlabel metal3 24024 15064 24024 15064 0 _0097_
rlabel metal3 29344 13944 29344 13944 0 _0098_
rlabel metal2 30520 14392 30520 14392 0 _0099_
rlabel metal2 31192 12544 31192 12544 0 _0100_
rlabel metal2 31640 14336 31640 14336 0 _0101_
rlabel metal2 30296 13160 30296 13160 0 _0102_
rlabel metal2 31248 13720 31248 13720 0 _0103_
rlabel metal3 30632 15064 30632 15064 0 _0104_
rlabel metal2 30688 13944 30688 13944 0 _0105_
rlabel metal2 29176 19320 29176 19320 0 _0106_
rlabel metal3 35000 21672 35000 21672 0 _0107_
rlabel metal3 31976 19992 31976 19992 0 _0108_
rlabel metal2 31528 21056 31528 21056 0 _0109_
rlabel metal2 31304 21616 31304 21616 0 _0110_
rlabel metal2 29792 20776 29792 20776 0 _0111_
rlabel metal2 26600 18928 26600 18928 0 _0112_
rlabel metal2 26992 17752 26992 17752 0 _0113_
rlabel metal2 29400 23856 29400 23856 0 _0114_
rlabel metal2 27664 20104 27664 20104 0 _0115_
rlabel metal2 18984 16352 18984 16352 0 _0116_
rlabel metal3 32704 26264 32704 26264 0 _0117_
rlabel metal3 34328 19992 34328 19992 0 _0118_
rlabel metal2 35056 19992 35056 19992 0 _0119_
rlabel metal2 34608 20216 34608 20216 0 _0120_
rlabel metal2 27160 7420 27160 7420 0 _0121_
rlabel metal2 23800 9184 23800 9184 0 _0122_
rlabel metal3 24696 9128 24696 9128 0 _0123_
rlabel metal2 20440 11760 20440 11760 0 _0124_
rlabel metal2 22344 9856 22344 9856 0 _0125_
rlabel metal2 25592 10248 25592 10248 0 _0126_
rlabel metal2 27608 8120 27608 8120 0 _0127_
rlabel metal2 24584 9912 24584 9912 0 _0128_
rlabel metal2 26040 9912 26040 9912 0 _0129_
rlabel metal2 25704 12320 25704 12320 0 _0130_
rlabel metal2 26908 13832 26908 13832 0 _0131_
rlabel metal2 27944 12768 27944 12768 0 _0132_
rlabel metal2 25368 14000 25368 14000 0 _0133_
rlabel metal3 24640 15176 24640 15176 0 _0134_
rlabel metal2 29176 11648 29176 11648 0 _0135_
rlabel metal3 28896 11256 28896 11256 0 _0136_
rlabel metal2 28112 8680 28112 8680 0 _0137_
rlabel metal2 32312 9128 32312 9128 0 _0138_
rlabel metal3 24864 9576 24864 9576 0 _0139_
rlabel metal2 24248 10192 24248 10192 0 _0140_
rlabel metal2 25200 9128 25200 9128 0 _0141_
rlabel metal2 26936 9520 26936 9520 0 _0142_
rlabel metal2 28448 8456 28448 8456 0 _0143_
rlabel metal3 28616 10696 28616 10696 0 _0144_
rlabel metal2 29512 10304 29512 10304 0 _0145_
rlabel metal2 29960 11648 29960 11648 0 _0146_
rlabel metal3 28224 14616 28224 14616 0 _0147_
rlabel metal2 27496 13608 27496 13608 0 _0148_
rlabel metal2 28168 11592 28168 11592 0 _0149_
rlabel metal2 28616 10864 28616 10864 0 _0150_
rlabel metal2 27832 9464 27832 9464 0 _0151_
rlabel metal2 27944 10080 27944 10080 0 _0152_
rlabel metal2 27608 12264 27608 12264 0 _0153_
rlabel metal3 28280 16296 28280 16296 0 _0154_
rlabel metal2 18704 9912 18704 9912 0 _0155_
rlabel metal2 25480 12600 25480 12600 0 _0156_
rlabel metal2 24360 11312 24360 11312 0 _0157_
rlabel metal3 25984 11928 25984 11928 0 _0158_
rlabel metal2 26712 13384 26712 13384 0 _0159_
rlabel metal3 28840 16968 28840 16968 0 _0160_
rlabel metal3 19152 23688 19152 23688 0 _0161_
rlabel metal2 18424 33264 18424 33264 0 _0162_
rlabel metal3 17416 33544 17416 33544 0 _0163_
rlabel metal2 19656 33684 19656 33684 0 _0164_
rlabel metal2 19096 32480 19096 32480 0 _0165_
rlabel metal3 18032 34216 18032 34216 0 _0166_
rlabel metal2 21448 31696 21448 31696 0 _0167_
rlabel metal2 23576 31808 23576 31808 0 _0168_
rlabel metal2 31976 29680 31976 29680 0 _0169_
rlabel metal2 32536 39088 32536 39088 0 _0170_
rlabel metal2 30968 38976 30968 38976 0 _0171_
rlabel metal2 33656 29680 33656 29680 0 _0172_
rlabel metal2 30576 29512 30576 29512 0 _0173_
rlabel metal2 31584 26264 31584 26264 0 _0174_
rlabel metal2 37016 30296 37016 30296 0 _0175_
rlabel metal3 37072 29400 37072 29400 0 _0176_
rlabel metal3 32480 30072 32480 30072 0 _0177_
rlabel metal2 23800 31248 23800 31248 0 _0178_
rlabel metal2 15176 37688 15176 37688 0 _0179_
rlabel metal2 15288 34552 15288 34552 0 _0180_
rlabel metal2 23240 32256 23240 32256 0 _0181_
rlabel metal2 21560 31584 21560 31584 0 _0182_
rlabel metal3 20664 23912 20664 23912 0 _0183_
rlabel metal3 16632 23688 16632 23688 0 _0184_
rlabel metal2 20216 24080 20216 24080 0 _0185_
rlabel metal3 23800 20776 23800 20776 0 _0186_
rlabel metal2 26040 19880 26040 19880 0 _0187_
rlabel metal2 31864 12488 31864 12488 0 _0188_
rlabel metal2 32144 19992 32144 19992 0 _0189_
rlabel metal2 33320 21056 33320 21056 0 _0190_
rlabel metal2 20216 18984 20216 18984 0 _0191_
rlabel metal3 19152 20104 19152 20104 0 _0192_
rlabel metal2 19712 11592 19712 11592 0 _0193_
rlabel metal2 19544 18424 19544 18424 0 _0194_
rlabel metal2 20328 19040 20328 19040 0 _0195_
rlabel metal3 19152 18536 19152 18536 0 _0196_
rlabel metal2 8904 22064 8904 22064 0 _0197_
rlabel metal2 10360 24752 10360 24752 0 _0198_
rlabel metal2 14616 8680 14616 8680 0 _0199_
rlabel metal3 17472 18424 17472 18424 0 _0200_
rlabel metal2 20776 19600 20776 19600 0 _0201_
rlabel metal2 23912 31248 23912 31248 0 _0202_
rlabel metal2 18872 9128 18872 9128 0 _0203_
rlabel metal3 19712 8344 19712 8344 0 _0204_
rlabel via2 21336 8232 21336 8232 0 _0205_
rlabel metal2 23128 5600 23128 5600 0 _0206_
rlabel metal2 26824 22064 26824 22064 0 _0207_
rlabel metal2 26376 22232 26376 22232 0 _0208_
rlabel metal2 21392 5320 21392 5320 0 _0209_
rlabel metal2 24136 4816 24136 4816 0 _0210_
rlabel metal2 24248 6160 24248 6160 0 _0211_
rlabel metal2 24416 4424 24416 4424 0 _0212_
rlabel metal2 24696 6384 24696 6384 0 _0213_
rlabel metal2 21896 23520 21896 23520 0 _0214_
rlabel metal2 5376 20104 5376 20104 0 _0215_
rlabel metal2 2408 20384 2408 20384 0 _0216_
rlabel metal2 3248 19432 3248 19432 0 _0217_
rlabel metal2 3080 20216 3080 20216 0 _0218_
rlabel metal2 4760 22288 4760 22288 0 _0219_
rlabel metal2 9072 22904 9072 22904 0 _0220_
rlabel metal2 10192 11256 10192 11256 0 _0221_
rlabel metal2 12208 9912 12208 9912 0 _0222_
rlabel metal3 15624 12376 15624 12376 0 _0223_
rlabel metal2 9856 15288 9856 15288 0 _0224_
rlabel metal2 8512 19992 8512 19992 0 _0225_
rlabel metal2 18536 24472 18536 24472 0 _0226_
rlabel metal2 9016 15456 9016 15456 0 _0227_
rlabel metal2 11256 12936 11256 12936 0 _0228_
rlabel metal2 7672 11088 7672 11088 0 _0229_
rlabel metal2 4088 18648 4088 18648 0 _0230_
rlabel metal2 2856 20328 2856 20328 0 _0231_
rlabel metal2 4536 18312 4536 18312 0 _0232_
rlabel metal3 6496 21784 6496 21784 0 _0233_
rlabel metal2 7896 12600 7896 12600 0 _0234_
rlabel metal4 6328 17360 6328 17360 0 _0235_
rlabel metal2 7560 11088 7560 11088 0 _0236_
rlabel metal2 9800 10864 9800 10864 0 _0237_
rlabel metal2 11592 12488 11592 12488 0 _0238_
rlabel metal2 9688 10864 9688 10864 0 _0239_
rlabel metal2 8792 12544 8792 12544 0 _0240_
rlabel metal2 22792 30072 22792 30072 0 _0241_
rlabel metal3 7168 23912 7168 23912 0 _0242_
rlabel metal2 7560 15792 7560 15792 0 _0243_
rlabel metal3 5768 15288 5768 15288 0 _0244_
rlabel metal3 8904 12040 8904 12040 0 _0245_
rlabel metal2 8456 12544 8456 12544 0 _0246_
rlabel metal2 6328 16240 6328 16240 0 _0247_
rlabel metal3 5320 14616 5320 14616 0 _0248_
rlabel metal2 5880 13440 5880 13440 0 _0249_
rlabel metal2 9688 13104 9688 13104 0 _0250_
rlabel metal3 8512 12712 8512 12712 0 _0251_
rlabel metal2 24360 27888 24360 27888 0 _0252_
rlabel metal2 8512 10584 8512 10584 0 _0253_
rlabel metal3 6776 16072 6776 16072 0 _0254_
rlabel metal3 6496 14504 6496 14504 0 _0255_
rlabel metal2 5768 14448 5768 14448 0 _0256_
rlabel metal2 6104 14280 6104 14280 0 _0257_
rlabel metal2 8456 14168 8456 14168 0 _0258_
rlabel metal2 8680 10808 8680 10808 0 _0259_
rlabel metal2 22568 27608 22568 27608 0 _0260_
rlabel metal2 3248 16856 3248 16856 0 _0261_
rlabel metal2 5768 16688 5768 16688 0 _0262_
rlabel metal2 7224 15232 7224 15232 0 _0263_
rlabel metal2 5992 18928 5992 18928 0 _0264_
rlabel metal2 7784 19208 7784 19208 0 _0265_
rlabel metal3 8064 15512 8064 15512 0 _0266_
rlabel metal3 8288 16856 8288 16856 0 _0267_
rlabel metal2 5656 16688 5656 16688 0 _0268_
rlabel metal2 6104 16856 6104 16856 0 _0269_
rlabel metal3 7728 18424 7728 18424 0 _0270_
rlabel metal2 7112 16464 7112 16464 0 _0271_
rlabel metal2 7896 16184 7896 16184 0 _0272_
rlabel metal2 7560 16408 7560 16408 0 _0273_
rlabel metal2 17528 35560 17528 35560 0 _0274_
rlabel metal3 6384 20776 6384 20776 0 _0275_
rlabel metal3 11032 19208 11032 19208 0 _0276_
rlabel metal2 6328 19040 6328 19040 0 _0277_
rlabel metal2 7448 18816 7448 18816 0 _0278_
rlabel metal2 7336 18704 7336 18704 0 _0279_
rlabel metal3 8120 18984 8120 18984 0 _0280_
rlabel metal2 7000 17864 7000 17864 0 _0281_
rlabel metal2 7224 17808 7224 17808 0 _0282_
rlabel metal2 8232 18816 8232 18816 0 _0283_
rlabel metal3 8680 19208 8680 19208 0 _0284_
rlabel metal2 9576 19824 9576 19824 0 _0285_
rlabel metal3 7448 23352 7448 23352 0 _0286_
rlabel metal2 6888 21952 6888 21952 0 _0287_
rlabel metal2 5656 20272 5656 20272 0 _0288_
rlabel metal2 6216 21280 6216 21280 0 _0289_
rlabel metal2 6776 21840 6776 21840 0 _0290_
rlabel metal3 6272 23240 6272 23240 0 _0291_
rlabel metal2 6328 22400 6328 22400 0 _0292_
rlabel metal2 6440 22512 6440 22512 0 _0293_
rlabel metal2 5320 23408 5320 23408 0 _0294_
rlabel metal2 22232 31360 22232 31360 0 _0295_
rlabel metal2 7112 24808 7112 24808 0 _0296_
rlabel metal2 4200 24360 4200 24360 0 _0297_
rlabel metal2 6608 23352 6608 23352 0 _0298_
rlabel metal2 5208 21280 5208 21280 0 _0299_
rlabel metal2 5880 19712 5880 19712 0 _0300_
rlabel metal2 5992 22400 5992 22400 0 _0301_
rlabel metal3 5040 23128 5040 23128 0 _0302_
rlabel metal2 4760 23520 4760 23520 0 _0303_
rlabel metal2 5656 22176 5656 22176 0 _0304_
rlabel metal2 6440 23464 6440 23464 0 _0305_
rlabel metal2 6776 23968 6776 23968 0 _0306_
rlabel metal2 6552 24976 6552 24976 0 _0307_
rlabel metal3 9240 29400 9240 29400 0 _0308_
rlabel metal2 16408 34608 16408 34608 0 _0309_
rlabel metal2 9744 28056 9744 28056 0 _0310_
rlabel metal3 25200 31752 25200 31752 0 _0311_
rlabel metal2 24696 31696 24696 31696 0 _0312_
rlabel metal2 8904 29792 8904 29792 0 _0313_
rlabel metal2 8064 29512 8064 29512 0 _0314_
rlabel metal2 5992 29568 5992 29568 0 _0315_
rlabel metal3 12936 37800 12936 37800 0 _0316_
rlabel metal2 15960 31976 15960 31976 0 _0317_
rlabel metal3 16632 33320 16632 33320 0 _0318_
rlabel metal2 10584 33376 10584 33376 0 _0319_
rlabel metal2 9576 30464 9576 30464 0 _0320_
rlabel metal3 9688 34048 9688 34048 0 _0321_
rlabel metal2 8624 32760 8624 32760 0 _0322_
rlabel metal3 8400 32424 8400 32424 0 _0323_
rlabel metal2 16184 27832 16184 27832 0 _0324_
rlabel metal3 16072 34104 16072 34104 0 _0325_
rlabel metal3 15288 37296 15288 37296 0 _0326_
rlabel metal2 13608 34496 13608 34496 0 _0327_
rlabel metal2 18984 35560 18984 35560 0 _0328_
rlabel metal2 11368 33600 11368 33600 0 _0329_
rlabel metal2 9856 34328 9856 34328 0 _0330_
rlabel metal2 9800 36008 9800 36008 0 _0331_
rlabel metal2 21896 36400 21896 36400 0 _0332_
rlabel metal3 11032 36568 11032 36568 0 _0333_
rlabel metal2 11816 34384 11816 34384 0 _0334_
rlabel metal2 11032 33768 11032 33768 0 _0335_
rlabel metal2 15624 37408 15624 37408 0 _0336_
rlabel metal2 15232 36568 15232 36568 0 _0337_
rlabel metal2 13720 36792 13720 36792 0 _0338_
rlabel metal3 13272 36568 13272 36568 0 _0339_
rlabel metal2 16352 37240 16352 37240 0 _0340_
rlabel metal2 16744 37576 16744 37576 0 _0341_
rlabel metal2 16184 37184 16184 37184 0 _0342_
rlabel metal2 16968 36680 16968 36680 0 _0343_
rlabel metal2 16632 36064 16632 36064 0 _0344_
rlabel metal2 16632 35448 16632 35448 0 _0345_
rlabel metal2 17360 35784 17360 35784 0 _0346_
rlabel metal2 15344 33432 15344 33432 0 _0347_
rlabel metal2 14672 34888 14672 34888 0 _0348_
rlabel metal2 15400 34552 15400 34552 0 _0349_
rlabel metal2 16296 34552 16296 34552 0 _0350_
rlabel metal2 14952 33824 14952 33824 0 _0351_
rlabel metal2 13832 33768 13832 33768 0 _0352_
rlabel metal2 25592 39144 25592 39144 0 _0353_
rlabel metal2 19544 34608 19544 34608 0 _0354_
rlabel metal2 19768 35224 19768 35224 0 _0355_
rlabel metal2 20888 36456 20888 36456 0 _0356_
rlabel metal2 21672 37184 21672 37184 0 _0357_
rlabel metal2 24136 28336 24136 28336 0 _0358_
rlabel metal2 24360 28728 24360 28728 0 _0359_
rlabel metal2 30856 40264 30856 40264 0 _0360_
rlabel metal2 26488 36736 26488 36736 0 _0361_
rlabel metal2 26376 37240 26376 37240 0 _0362_
rlabel metal2 24920 37184 24920 37184 0 _0363_
rlabel metal2 25200 38696 25200 38696 0 _0364_
rlabel metal2 31136 37240 31136 37240 0 _0365_
rlabel metal2 30184 39088 30184 39088 0 _0366_
rlabel metal2 27048 36960 27048 36960 0 _0367_
rlabel metal2 29960 39032 29960 39032 0 _0368_
rlabel metal2 28616 38696 28616 38696 0 _0369_
rlabel metal2 30352 40936 30352 40936 0 _0370_
rlabel metal2 27832 39480 27832 39480 0 _0371_
rlabel metal3 31416 37800 31416 37800 0 _0372_
rlabel metal3 33824 31752 33824 31752 0 _0373_
rlabel metal2 32200 32928 32200 32928 0 _0374_
rlabel metal2 30576 37464 30576 37464 0 _0375_
rlabel metal2 30072 39088 30072 39088 0 _0376_
rlabel metal2 29848 39200 29848 39200 0 _0377_
rlabel metal2 31528 39704 31528 39704 0 _0378_
rlabel metal3 30800 34328 30800 34328 0 _0379_
rlabel metal3 32480 38696 32480 38696 0 _0380_
rlabel metal2 31192 37464 31192 37464 0 _0381_
rlabel metal3 31696 35784 31696 35784 0 _0382_
rlabel metal3 30072 33320 30072 33320 0 _0383_
rlabel metal2 33152 34216 33152 34216 0 _0384_
rlabel metal3 32816 35672 32816 35672 0 _0385_
rlabel metal2 32200 35504 32200 35504 0 _0386_
rlabel metal2 30856 35168 30856 35168 0 _0387_
rlabel metal2 31416 34440 31416 34440 0 _0388_
rlabel metal2 31528 32088 31528 32088 0 _0389_
rlabel metal3 31304 33544 31304 33544 0 _0390_
rlabel metal2 31192 33040 31192 33040 0 _0391_
rlabel metal2 29512 32872 29512 32872 0 _0392_
rlabel metal3 27440 32536 27440 32536 0 _0393_
rlabel metal2 24584 31472 24584 31472 0 _0394_
rlabel metal2 25592 32480 25592 32480 0 _0395_
rlabel metal2 25592 18424 25592 18424 0 _0396_
rlabel metal2 35336 31584 35336 31584 0 _0397_
rlabel metal2 31192 32536 31192 32536 0 _0398_
rlabel metal3 35560 33208 35560 33208 0 _0399_
rlabel metal2 37072 32760 37072 32760 0 _0400_
rlabel metal2 37800 32872 37800 32872 0 _0401_
rlabel metal2 37520 32536 37520 32536 0 _0402_
rlabel metal3 37464 31864 37464 31864 0 _0403_
rlabel metal2 30520 23240 30520 23240 0 _0404_
rlabel metal2 36680 30352 36680 30352 0 _0405_
rlabel metal2 36568 31416 36568 31416 0 _0406_
rlabel metal2 36008 32144 36008 32144 0 _0407_
rlabel metal3 34832 32424 34832 32424 0 _0408_
rlabel metal2 35560 31808 35560 31808 0 _0409_
rlabel metal2 37688 30632 37688 30632 0 _0410_
rlabel metal2 26712 29288 26712 29288 0 _0411_
rlabel metal2 33600 31752 33600 31752 0 _0412_
rlabel metal2 28056 30856 28056 30856 0 _0413_
rlabel metal2 27832 31136 27832 31136 0 _0414_
rlabel metal2 27496 31024 27496 31024 0 _0415_
rlabel metal2 26600 31192 26600 31192 0 _0416_
rlabel metal2 26824 30576 26824 30576 0 _0417_
rlabel metal2 25928 30464 25928 30464 0 _0418_
rlabel metal3 23688 23912 23688 23912 0 _0419_
rlabel metal2 24472 23520 24472 23520 0 _0420_
rlabel metal2 21448 14728 21448 14728 0 _0421_
rlabel metal2 15288 12992 15288 12992 0 _0422_
rlabel metal2 13720 12824 13720 12824 0 _0423_
rlabel metal2 12488 14784 12488 14784 0 _0424_
rlabel metal3 13216 14504 13216 14504 0 _0425_
rlabel metal2 13496 11984 13496 11984 0 _0426_
rlabel metal2 15624 14112 15624 14112 0 _0427_
rlabel metal3 15120 13608 15120 13608 0 _0428_
rlabel metal2 15512 14224 15512 14224 0 _0429_
rlabel metal3 14448 14392 14448 14392 0 _0430_
rlabel metal2 14168 18200 14168 18200 0 _0431_
rlabel metal2 14504 19376 14504 19376 0 _0432_
rlabel metal2 12096 20104 12096 20104 0 _0433_
rlabel metal3 13496 20104 13496 20104 0 _0434_
rlabel metal2 15400 22008 15400 22008 0 _0435_
rlabel metal2 12824 20272 12824 20272 0 _0436_
rlabel metal2 13608 19992 13608 19992 0 _0437_
rlabel metal2 15064 19488 15064 19488 0 _0438_
rlabel metal3 19880 19208 19880 19208 0 _0439_
rlabel metal2 32984 25648 32984 25648 0 _0440_
rlabel metal2 33040 26376 33040 26376 0 _0441_
rlabel metal2 33040 29400 33040 29400 0 _0442_
rlabel metal2 33320 24920 33320 24920 0 _0443_
rlabel metal2 36344 26600 36344 26600 0 _0444_
rlabel metal3 32200 24696 32200 24696 0 _0445_
rlabel metal2 33544 25480 33544 25480 0 _0446_
rlabel metal2 32256 24808 32256 24808 0 _0447_
rlabel metal2 32312 26376 32312 26376 0 _0448_
rlabel metal2 31472 26488 31472 26488 0 _0449_
rlabel metal2 35840 27832 35840 27832 0 _0450_
rlabel metal2 36344 27496 36344 27496 0 _0451_
rlabel metal2 32032 27272 32032 27272 0 _0452_
rlabel metal2 28056 27328 28056 27328 0 _0453_
rlabel metal2 26712 27384 26712 27384 0 _0454_
rlabel metal3 29848 27944 29848 27944 0 _0455_
rlabel metal2 33096 27160 33096 27160 0 _0456_
rlabel metal2 36008 28168 36008 28168 0 _0457_
rlabel metal2 34888 26628 34888 26628 0 _0458_
rlabel metal2 33544 27552 33544 27552 0 _0459_
rlabel metal2 32200 27440 32200 27440 0 _0460_
rlabel metal2 30072 27104 30072 27104 0 _0461_
rlabel metal2 34608 25592 34608 25592 0 _0462_
rlabel metal2 33880 27552 33880 27552 0 _0463_
rlabel metal2 31864 26376 31864 26376 0 _0464_
rlabel metal2 29848 27384 29848 27384 0 _0465_
rlabel metal2 29512 29568 29512 29568 0 _0466_
rlabel metal2 29512 28112 29512 28112 0 _0467_
rlabel metal3 18816 26488 18816 26488 0 _0468_
rlabel metal2 18312 27104 18312 27104 0 _0469_
rlabel metal3 17752 26880 17752 26880 0 _0470_
rlabel metal2 28952 22512 28952 22512 0 _0471_
rlabel metal2 27832 22680 27832 22680 0 _0472_
rlabel metal2 19768 26488 19768 26488 0 _0473_
rlabel metal2 17752 28112 17752 28112 0 _0474_
rlabel metal2 15736 29008 15736 29008 0 _0475_
rlabel metal2 19880 29008 19880 29008 0 _0476_
rlabel metal2 12936 27776 12936 27776 0 _0477_
rlabel metal3 12768 28504 12768 28504 0 _0478_
rlabel metal2 18088 29176 18088 29176 0 _0479_
rlabel metal3 18648 32536 18648 32536 0 _0480_
rlabel metal3 17584 31752 17584 31752 0 _0481_
rlabel metal3 17360 30184 17360 30184 0 _0482_
rlabel metal2 18088 28784 18088 28784 0 _0483_
rlabel metal2 19432 29288 19432 29288 0 _0484_
rlabel metal2 19712 27048 19712 27048 0 _0485_
rlabel metal3 20048 27048 20048 27048 0 _0486_
rlabel metal2 18648 32200 18648 32200 0 _0487_
rlabel metal2 20776 30688 20776 30688 0 _0488_
rlabel metal3 20944 29400 20944 29400 0 _0489_
rlabel metal2 20888 29456 20888 29456 0 _0490_
rlabel metal2 16800 27048 16800 27048 0 _0491_
rlabel metal2 18984 28560 18984 28560 0 _0492_
rlabel metal2 19152 31192 19152 31192 0 _0493_
rlabel metal2 19264 30968 19264 30968 0 _0494_
rlabel metal2 18312 30072 18312 30072 0 _0495_
rlabel metal2 17640 27888 17640 27888 0 _0496_
rlabel metal2 16688 29176 16688 29176 0 _0497_
rlabel metal2 18592 29400 18592 29400 0 _0498_
rlabel metal2 19152 29624 19152 29624 0 _0499_
rlabel metal2 20216 27720 20216 27720 0 _0500_
rlabel metal2 31752 12040 31752 12040 0 _0501_
rlabel metal3 33544 21336 33544 21336 0 _0502_
rlabel metal2 34776 9744 34776 9744 0 _0503_
rlabel metal3 33936 9688 33936 9688 0 _0504_
rlabel metal3 33208 13160 33208 13160 0 _0505_
rlabel metal2 32312 14112 32312 14112 0 _0506_
rlabel metal3 31864 12936 31864 12936 0 _0507_
rlabel metal2 33768 13636 33768 13636 0 _0508_
rlabel metal2 33656 13104 33656 13104 0 _0509_
rlabel metal3 35168 16856 35168 16856 0 _0510_
rlabel metal2 34272 16296 34272 16296 0 _0511_
rlabel metal2 36568 17248 36568 17248 0 _0512_
rlabel metal3 35616 18312 35616 18312 0 _0513_
rlabel metal2 36120 18144 36120 18144 0 _0514_
rlabel metal2 37240 21616 37240 21616 0 _0515_
rlabel metal2 37016 21616 37016 21616 0 _0516_
rlabel metal2 37856 19432 37856 19432 0 _0517_
rlabel metal2 38248 22400 38248 22400 0 _0518_
rlabel metal2 38024 22176 38024 22176 0 _0519_
rlabel metal2 11760 20104 11760 20104 0 _0520_
rlabel metal2 10808 19656 10808 19656 0 _0521_
rlabel metal2 11144 19712 11144 19712 0 _0522_
rlabel metal3 13440 19992 13440 19992 0 _0523_
rlabel metal2 12040 19656 12040 19656 0 _0524_
rlabel metal3 13384 18424 13384 18424 0 _0525_
rlabel metal2 24920 18648 24920 18648 0 _0526_
rlabel metal3 25088 18424 25088 18424 0 _0527_
rlabel metal3 17360 11368 17360 11368 0 _0528_
rlabel metal2 19320 12376 19320 12376 0 _0529_
rlabel metal3 17080 11592 17080 11592 0 _0530_
rlabel metal2 21336 22736 21336 22736 0 _0531_
rlabel metal2 19656 12488 19656 12488 0 _0532_
rlabel metal2 20552 12432 20552 12432 0 _0533_
rlabel metal3 18984 12936 18984 12936 0 _0534_
rlabel metal2 17192 11760 17192 11760 0 _0535_
rlabel metal2 19096 13888 19096 13888 0 _0536_
rlabel metal3 18648 12152 18648 12152 0 _0537_
rlabel metal3 17416 16296 17416 16296 0 _0538_
rlabel metal3 19376 15288 19376 15288 0 _0539_
rlabel metal2 19432 14616 19432 14616 0 _0540_
rlabel metal3 20944 15512 20944 15512 0 _0541_
rlabel metal2 16576 17080 16576 17080 0 _0542_
rlabel metal2 17360 19096 17360 19096 0 _0543_
rlabel metal2 17808 23912 17808 23912 0 _0544_
rlabel metal2 18088 24360 18088 24360 0 _0545_
rlabel metal2 17752 23184 17752 23184 0 _0546_
rlabel metal2 15736 22512 15736 22512 0 _0547_
rlabel metal2 15960 22680 15960 22680 0 _0548_
rlabel metal2 21560 21224 21560 21224 0 _0549_
rlabel metal2 20664 20272 20664 20272 0 _0550_
rlabel metal2 21840 19992 21840 19992 0 _0551_
rlabel metal2 21448 19656 21448 19656 0 _0552_
rlabel metal3 39634 14840 39634 14840 0 blue
rlabel metal2 31192 14560 31192 14560 0 clknet_0_wb_clk_i
rlabel metal2 19544 4704 19544 4704 0 clknet_3_0__leaf_wb_clk_i
rlabel metal2 2408 10528 2408 10528 0 clknet_3_1__leaf_wb_clk_i
rlabel metal2 32704 8008 32704 8008 0 clknet_3_2__leaf_wb_clk_i
rlabel metal2 21560 17640 21560 17640 0 clknet_3_3__leaf_wb_clk_i
rlabel metal2 4760 25480 4760 25480 0 clknet_3_4__leaf_wb_clk_i
rlabel metal2 11424 38808 11424 38808 0 clknet_3_5__leaf_wb_clk_i
rlabel metal2 25256 28672 25256 28672 0 clknet_3_6__leaf_wb_clk_i
rlabel metal3 25200 39368 25200 39368 0 clknet_3_7__leaf_wb_clk_i
rlabel metal3 40586 12824 40586 12824 0 debug_design_reset
rlabel metal2 40040 7784 40040 7784 0 debug_gpio_ready
rlabel metal2 1736 20440 1736 20440 0 down_key_n
rlabel metal2 40040 26656 40040 26656 0 ext_reset_n
rlabel metal2 40152 5656 40152 5656 0 gpio_ready
rlabel metal2 40040 21168 40040 21168 0 green
rlabel metal3 40418 20216 40418 20216 0 hsync
rlabel metal2 39592 15064 39592 15064 0 io_oeb[13]
rlabel metal2 39704 16912 39704 16912 0 io_oeb[14]
rlabel metal3 39634 18200 39634 18200 0 io_oeb[15]
rlabel metal2 39760 15512 39760 15512 0 io_oeb[16]
rlabel metal2 39704 18648 39704 18648 0 io_oeb[17]
rlabel metal3 39746 16184 39746 16184 0 io_oeb[18]
rlabel metal2 2072 19992 2072 19992 0 net1
rlabel metal2 38696 6608 38696 6608 0 net10
rlabel metal2 39144 20664 39144 20664 0 net11
rlabel metal2 33432 20160 33432 20160 0 net12
rlabel metal2 38920 14784 38920 14784 0 net13
rlabel metal2 38920 16184 38920 16184 0 net14
rlabel metal2 29848 18816 29848 18816 0 net15
rlabel metal2 32872 16128 32872 16128 0 net16
rlabel metal3 38780 18424 38780 18424 0 net17
rlabel metal2 30856 16520 30856 16520 0 net18
rlabel metal3 28056 17528 28056 17528 0 net19
rlabel metal2 39816 26712 39816 26712 0 net2
rlabel metal2 2968 24024 2968 24024 0 net20
rlabel metal3 20048 3528 20048 3528 0 net21
rlabel metal3 29344 17640 29344 17640 0 net22
rlabel metal2 29960 16912 29960 16912 0 net23
rlabel metal3 30856 17528 30856 17528 0 net24
rlabel metal3 30408 13608 30408 13608 0 net25
rlabel metal3 38920 12992 38920 12992 0 net26
rlabel metal3 26152 30184 26152 30184 0 net27
rlabel metal2 40152 37184 40152 37184 0 net28
rlabel metal2 32984 2030 32984 2030 0 net29
rlabel metal2 38472 5544 38472 5544 0 net3
rlabel metal3 40418 41048 40418 41048 0 net30
rlabel metal2 35672 44198 35672 44198 0 net31
rlabel metal2 10808 2030 10808 2030 0 net32
rlabel metal3 1246 5432 1246 5432 0 net33
rlabel metal2 40152 4816 40152 4816 0 net34
rlabel metal2 40152 4256 40152 4256 0 net35
rlabel metal2 10136 2030 10136 2030 0 net36
rlabel metal2 39256 2688 39256 2688 0 net37
rlabel metal3 854 6104 854 6104 0 net38
rlabel metal2 1736 3360 1736 3360 0 net39
rlabel metal2 2072 25872 2072 25872 0 net4
rlabel metal2 40208 40936 40208 40936 0 net40
rlabel metal2 40152 12208 40152 12208 0 net41
rlabel metal2 40152 42280 40152 42280 0 net42
rlabel metal2 40152 7896 40152 7896 0 net43
rlabel metal2 40152 40096 40152 40096 0 net44
rlabel metal2 39704 3584 39704 3584 0 net45
rlabel metal2 8120 44198 8120 44198 0 net46
rlabel metal3 1246 36344 1246 36344 0 net47
rlabel metal3 1246 4760 1246 4760 0 net48
rlabel metal2 40152 38640 40152 38640 0 net49
rlabel metal2 19992 19152 19992 19152 0 net5
rlabel metal2 40152 6272 40152 6272 0 net50
rlabel metal3 1246 40376 1246 40376 0 net51
rlabel metal2 40152 37744 40152 37744 0 net52
rlabel metal2 39256 41888 39256 41888 0 net53
rlabel metal3 1246 37016 1246 37016 0 net54
rlabel metal2 40208 39368 40208 39368 0 net55
rlabel metal2 38808 42616 38808 42616 0 net56
rlabel metal3 1246 4088 1246 4088 0 net57
rlabel metal2 39704 7168 39704 7168 0 net58
rlabel metal3 40152 3360 40152 3360 0 net59
rlabel metal2 3024 19320 3024 19320 0 net6
rlabel metal2 39816 25816 39816 25816 0 net7
rlabel metal2 29512 16408 29512 16408 0 net8
rlabel metal3 23968 24808 23968 24808 0 net9
rlabel metal2 1848 25592 1848 25592 0 new_game_n
rlabel metal3 19936 3416 19936 3416 0 pause_n
rlabel metal2 40040 19432 40040 19432 0 red
rlabel metal2 29568 23016 29568 23016 0 solo_squash.ballDirX
rlabel metal2 11480 31304 11480 31304 0 solo_squash.ballDirY
rlabel metal2 26656 34888 26656 34888 0 solo_squash.ballX\[0\]
rlabel metal2 26264 39704 26264 39704 0 solo_squash.ballX\[1\]
rlabel metal2 28728 39928 28728 39928 0 solo_squash.ballX\[2\]
rlabel metal2 32760 39928 32760 39928 0 solo_squash.ballX\[3\]
rlabel metal2 33992 34552 33992 34552 0 solo_squash.ballX\[4\]
rlabel metal2 29288 30016 29288 30016 0 solo_squash.ballX\[5\]
rlabel metal2 40152 30576 40152 30576 0 solo_squash.ballX\[6\]
rlabel metal2 38584 28952 38584 28952 0 solo_squash.ballX\[7\]
rlabel metal3 31808 26152 31808 26152 0 solo_squash.ballX\[8\]
rlabel metal3 10920 28728 10920 28728 0 solo_squash.ballY\[0\]
rlabel metal2 10472 28840 10472 28840 0 solo_squash.ballY\[1\]
rlabel metal2 8792 33768 8792 33768 0 solo_squash.ballY\[2\]
rlabel metal2 10808 35728 10808 35728 0 solo_squash.ballY\[3\]
rlabel metal2 14224 38696 14224 38696 0 solo_squash.ballY\[4\]
rlabel metal3 16968 36456 16968 36456 0 solo_squash.ballY\[5\]
rlabel metal3 15512 31864 15512 31864 0 solo_squash.ballY\[6\]
rlabel metal2 20496 35672 20496 35672 0 solo_squash.ballY\[7\]
rlabel metal2 30968 11816 30968 11816 0 solo_squash.h\[0\]
rlabel metal2 33096 9240 33096 9240 0 solo_squash.h\[1\]
rlabel metal2 28112 8232 28112 8232 0 solo_squash.h\[2\]
rlabel metal2 29904 12712 29904 12712 0 solo_squash.h\[3\]
rlabel metal2 29848 14616 29848 14616 0 solo_squash.h\[4\]
rlabel metal2 40152 16632 40152 16632 0 solo_squash.h\[5\]
rlabel metal2 40040 17360 40040 17360 0 solo_squash.h\[6\]
rlabel metal3 33376 20776 33376 20776 0 solo_squash.h\[7\]
rlabel metal2 40152 21224 40152 21224 0 solo_squash.h\[8\]
rlabel metal2 35784 25424 35784 25424 0 solo_squash.h\[9\]
rlabel metal3 21504 23800 21504 23800 0 solo_squash.hit
rlabel metal3 30576 25480 30576 25480 0 solo_squash.inBallX
rlabel metal3 20328 27160 20328 27160 0 solo_squash.inBallY
rlabel metal2 24696 19376 24696 19376 0 solo_squash.inPaddle
rlabel metal2 19320 8568 19320 8568 0 solo_squash.offset\[0\]
rlabel metal2 22456 7896 22456 7896 0 solo_squash.offset\[1\]
rlabel metal2 22344 8120 22344 8120 0 solo_squash.offset\[2\]
rlabel metal2 26040 6328 26040 6328 0 solo_squash.offset\[3\]
rlabel metal2 27496 6776 27496 6776 0 solo_squash.offset\[4\]
rlabel metal2 12936 10976 12936 10976 0 solo_squash.paddle\[0\]
rlabel metal3 5208 12936 5208 12936 0 solo_squash.paddle\[1\]
rlabel metal2 5152 10472 5152 10472 0 solo_squash.paddle\[2\]
rlabel metal2 6328 12432 6328 12432 0 solo_squash.paddle\[3\]
rlabel metal2 10360 13664 10360 13664 0 solo_squash.paddle\[4\]
rlabel metal2 4424 17192 4424 17192 0 solo_squash.paddle\[5\]
rlabel metal2 13608 19488 13608 19488 0 solo_squash.paddle\[6\]
rlabel metal3 2408 21784 2408 21784 0 solo_squash.paddle\[7\]
rlabel metal2 1736 25368 1736 25368 0 solo_squash.paddle\[8\]
rlabel metal3 20216 9688 20216 9688 0 solo_squash.v\[0\]
rlabel metal3 21168 9912 21168 9912 0 solo_squash.v\[1\]
rlabel metal3 20664 9576 20664 9576 0 solo_squash.v\[2\]
rlabel metal3 25088 13944 25088 13944 0 solo_squash.v\[3\]
rlabel metal2 13384 15232 13384 15232 0 solo_squash.v\[4\]
rlabel metal2 16072 19152 16072 19152 0 solo_squash.v\[5\]
rlabel metal2 16632 24752 16632 24752 0 solo_squash.v\[6\]
rlabel metal2 15848 22624 15848 22624 0 solo_squash.v\[7\]
rlabel metal3 20104 22344 20104 22344 0 solo_squash.v\[8\]
rlabel metal2 19488 17528 19488 17528 0 solo_squash.v\[9\]
rlabel metal2 1960 24136 1960 24136 0 speaker
rlabel metal2 1736 19376 1736 19376 0 up_key_n
rlabel metal3 20384 3640 20384 3640 0 vsync
rlabel metal3 2534 39704 2534 39704 0 wb_clk_i
rlabel metal2 40152 26600 40152 26600 0 wb_rst_i
<< properties >>
string FIXED_BBOX 0 0 41901 45485
<< end >>
